module debug(A_0_0, B_0_0, S_0_0, A_0_1, B_0_1, S_0_1, A_0_2, B_0_2, S_0_2, A_1_0, B_1_0, S_1_0, A_1_1, B_1_1, S_1_1, A_1_2, B_1_2, S_1_2, A_2_0, B_2_0, S_2_0, A_2_1, B_2_1, S_2_1, A_2_2, B_2_2, S_2_2, Cin_0, Cin_1, Cin_2, Cout_0, Cout_1, Cout_2);

   input A_0_0, A_0_1, A_0_2, A_1_0, A_1_1, A_1_2, A_2_0, A_2_1, A_2_2;
   input B_0_0, B_0_1, B_0_2, B_1_0, B_1_1, B_1_2, B_2_0, B_2_1, B_2_2;
   output S_0_0, S_0_1, S_0_2, S_1_0, S_1_1, S_1_2, S_2_0, S_2_1, S_2_2;
   input Cin_0, Cin_1, Cin_2;
   output Cout_0, Cout_1, Cout_2;
   wire W_0_0_1, W_0_0_2, W_0_0_3, W_0_0_4, W_0_1_1, W_0_1_2, W_0_1_3, W_0_1_4, W_0_2_1, W_0_2_2, W_0_2_3, W_0_2_4, W_1_0_1, W_1_0_2, W_1_0_3, W_1_0_4, W_1_1_1, W_1_1_2, W_1_1_3, W_1_1_4, W_1_2_1, W_1_2_2, W_1_2_3, W_1_2_4, W_2_0_1, W_2_0_2, W_2_0_3, W_2_0_4, W_2_1_1, W_2_1_2, W_2_1_3, W_2_1_4, W_2_2_1, W_2_2_2, W_2_2_3, W_2_2_4;
   GTECH_XOR2 u_0_0_1 (.A(A_0_0), .B(B_0_0), .Z(W_0_0_1));
   GTECH_XOR2 u_0_1_1 (.A(A_0_1), .B(B_0_1), .Z(W_0_1_1));
   GTECH_XOR2 u_0_2_1 (.A(A_0_2), .B(B_0_2), .Z(W_0_2_1));
   GTECH_XOR2 u_1_0_1 (.A(A_1_0), .B(B_1_0), .Z(W_1_0_1));
   GTECH_XOR2 u_1_1_1 (.A(A_1_1), .B(B_1_1), .Z(W_1_1_1));
   GTECH_XOR2 u_1_2_1 (.A(A_1_2), .B(B_1_2), .Z(W_1_2_1));
   GTECH_XOR2 u_2_0_1 (.A(A_2_0), .B(B_2_0), .Z(W_2_0_1));
   GTECH_XOR2 u_2_1_1 (.A(A_2_1), .B(B_2_1), .Z(W_2_1_1));
   GTECH_XOR2 u_2_2_1 (.A(A_2_2), .B(B_2_2), .Z(W_2_2_1));
   GTECH_AND2 u_0_0_2 (.A(A_0_0), .B(B_0_0), .Z(W_0_0_2));
   GTECH_AND2 u_0_1_2 (.A(A_0_1), .B(B_0_1), .Z(W_0_1_2));
   GTECH_AND2 u_0_2_2 (.A(A_0_2), .B(B_0_2), .Z(W_0_2_2));
   GTECH_AND2 u_1_0_2 (.A(A_1_0), .B(B_1_0), .Z(W_1_0_2));
   GTECH_AND2 u_1_1_2 (.A(A_1_1), .B(B_1_1), .Z(W_1_1_2));
   GTECH_AND2 u_1_2_2 (.A(A_1_2), .B(B_1_2), .Z(W_1_2_2));
   GTECH_AND2 u_2_0_2 (.A(A_2_0), .B(B_2_0), .Z(W_2_0_2));
   GTECH_AND2 u_2_1_2 (.A(A_2_1), .B(B_2_1), .Z(W_2_1_2));
   GTECH_AND2 u_2_2_2 (.A(A_2_2), .B(B_2_2), .Z(W_2_2_2));
   GTECH_AND2 u_0_0_3 (.A(W_0_0_1), .B(Cin_0), .Z(W_0_0_3));
   GTECH_AND2 u_0_1_3 (.A(W_0_1_1), .B(W_0_1_4), .Z(W_0_1_3));
   GTECH_AND2 u_0_2_3 (.A(W_0_2_1), .B(W_0_2_4), .Z(W_0_2_3));
   GTECH_AND2 u_1_0_3 (.A(W_1_0_1), .B(Cin_1), .Z(W_1_0_3));
   GTECH_AND2 u_1_1_3 (.A(W_1_1_1), .B(W_1_1_4), .Z(W_1_1_3));
   GTECH_AND2 u_1_2_3 (.A(W_1_2_1), .B(W_1_2_4), .Z(W_1_2_3));
   GTECH_AND2 u_2_0_3 (.A(W_2_0_1), .B(Cin_2), .Z(W_2_0_3));
   GTECH_AND2 u_2_1_3 (.A(W_2_1_1), .B(W_2_1_4), .Z(W_2_1_3));
   GTECH_AND2 u_2_2_3 (.A(W_2_2_1), .B(W_2_2_4), .Z(W_2_2_3));
   GTECH_XOR2 u_0_0_4 (.A(Cin_0), .B(W_0_0_1), .Z(S_0_0));
   GTECH_XOR2 u_0_1_4 (.A(W_0_1_4), .B(W_0_1_1), .Z(S_0_1));
   GTECH_XOR2 u_0_2_4 (.A(W_0_2_4), .B(W_0_2_1), .Z(S_0_2));
   GTECH_XOR2 u_1_0_4 (.A(Cin_1), .B(W_1_0_1), .Z(S_1_0));
   GTECH_XOR2 u_1_1_4 (.A(W_1_1_4), .B(W_1_1_1), .Z(S_1_1));
   GTECH_XOR2 u_1_2_4 (.A(W_1_2_4), .B(W_1_2_1), .Z(S_1_2));
   GTECH_XOR2 u_2_0_4 (.A(Cin_2), .B(W_2_0_1), .Z(S_2_0));
   GTECH_XOR2 u_2_1_4 (.A(W_2_1_4), .B(W_2_1_1), .Z(S_2_1));
   GTECH_XOR2 u_2_2_4 (.A(W_2_2_4), .B(W_2_2_1), .Z(S_2_2));
   GTECH_AND2 u_0_0_5 (.A(W_0_0_2), .B(W_0_0_3), .Z(W_0_1_4));
   GTECH_AND2 u_0_1_5 (.A(W_0_1_2), .B(W_0_1_3), .Z(W_0_2_4));
   GTECH_AND2 u_0_2_5 (.A(W_0_2_2), .B(W_0_2_3), .Z(Cout_0));
   GTECH_AND2 u_1_0_5 (.A(W_1_0_2), .B(W_1_0_3), .Z(W_1_1_4));
   GTECH_AND2 u_1_1_5 (.A(W_1_1_2), .B(W_1_1_3), .Z(W_1_2_4));
   GTECH_AND2 u_1_2_5 (.A(W_1_2_2), .B(W_1_2_3), .Z(Cout_1));
   GTECH_AND2 u_2_0_5 (.A(W_2_0_2), .B(W_2_0_3), .Z(W_2_1_4));
   GTECH_AND2 u_2_1_5 (.A(W_2_1_2), .B(W_2_1_3), .Z(W_2_2_4));
   GTECH_AND2 u_2_2_5 (.A(W_2_2_2), .B(W_2_2_3), .Z(Cout_2));

endmodule
