
module sec_1dDCT_seq_width8 ( x0, x1, x2, x3, x4, x5, x6, x7, clk, D0, D1, D2, 
        D3, D4, D5, D6, D7 );
  input [8:0] x0;
  input [8:0] x1;
  input [8:0] x2;
  input [8:0] x3;
  input [8:0] x4;
  input [8:0] x5;
  input [8:0] x6;
  input [8:0] x7;
  output [12:0] D0;
  output [12:0] D1;
  output [12:0] D2;
  output [12:0] D3;
  output [12:0] D4;
  output [12:0] D5;
  output [12:0] D6;
  output [12:0] D7;
  input clk;
  wire   \temp5t[0] , \temp6t[0] , \temp7t[0] , \temp8t[0] , \s6[0] , \s7[0] ,
         \U1/Ytt[11] , \U1/Ytt[10] , \U1/Ytt[9] , \U1/Ytt[8] , \U1/Ytt[7] ,
         \U1/Ytt[6] , \U1/Ytt[5] , \U1/Ytt[4] , \U1/Ytt[3] , \U1/Ytt[2] ,
         \U1/Ytt[1] , \U1/Ytt[0] , \U1/Xtt[11] , \U1/Xtt[10] , \U1/Xtt[9] ,
         \U1/Xtt[8] , \U1/Xtt[7] , \U1/Xtt[6] , \U1/Xtt[5] , \U1/Xtt[4] ,
         \U1/Xtt[3] , \U1/Xtt[2] , \U1/Xtt[1] , \U1/Xtt[0] , \U1/result6[13] ,
         \U1/result6[2] , \U1/result6[1] , \U1/result6[0] , \U1/result5[13] ,
         \U1/result5[2] , \U1/result5[1] , \U1/result5[0] , \U1/temp_yyyt[0] ,
         \U1/temp_yyyt[1] , \U1/temp_yyyt[2] , \U1/temp_yyyt[3] ,
         \U1/temp_yyyt[4] , \U1/temp_yyyt[5] , \U1/temp_yyyt[6] ,
         \U1/temp_yyyt[7] , \U1/temp_xxxt[0] , \U1/temp_xxxt[1] ,
         \U1/temp_xxxt[2] , \U1/temp_xxxt[3] , \U1/temp_xxxt[4] ,
         \U1/temp_xxxt[5] , \U1/temp_xxxt[6] , \U1/temp_xxxt[7] ,
         \U1/temp_yyy[11] , \U1/temp_yyy[10] , \U1/temp_yyy[9] ,
         \U1/temp_yyy[8] , \U1/temp_yyy[7] , \U1/temp_yyy[6] ,
         \U1/temp_yyy[5] , \U1/temp_yyy[4] , \U1/temp_yyy[3] ,
         \U1/temp_yyy[2] , \U1/temp_yyy[1] , \U1/temp_xxx[11] ,
         \U1/temp_xxx[10] , \U1/temp_xxx[9] , \U1/temp_xxx[8] ,
         \U1/temp_xxx[7] , \U1/temp_xxx[6] , \U1/temp_xxx[5] ,
         \U1/temp_xxx[4] , \U1/temp_xxx[3] , \U1/temp_xxx[2] ,
         \U1/temp_xxx[1] , \U1/temp_xxx[0] , \U2/Ytt[10] , \U2/Ytt[9] ,
         \U2/Ytt[8] , \U2/Ytt[7] , \U2/Ytt[6] , \U2/Ytt[5] , \U2/Ytt[4] ,
         \U2/Ytt[3] , \U2/Ytt[2] , \U2/Ytt[1] , \U2/Ytt[0] , \U2/Xtt[10] ,
         \U2/Xtt[9] , \U2/Xtt[8] , \U2/Xtt[7] , \U2/Xtt[6] , \U2/Xtt[5] ,
         \U2/Xtt[4] , \U2/Xtt[3] , \U2/Xtt[2] , \U2/Xtt[1] , \U2/Xtt[0] ,
         \U2/result2[11] , \U2/result2[9] , \U2/result2[8] , \U2/result2[7] ,
         \U2/result2[6] , \U2/result2[5] , \U2/result2[4] , \U2/result2[3] ,
         \U2/result2[2] , \U2/result2[1] , \U2/result2[0] , \U2/result1[11] ,
         \U2/result1[9] , \U2/result1[8] , \U2/result1[7] , \U2/result1[6] ,
         \U2/result1[5] , \U2/result1[4] , \U2/result1[3] , \U2/result1[2] ,
         \U2/result1[1] , \U2/result1[0] , \U2/temp_yt[0] , \U2/temp_xt[0] ,
         \U2/temp_y[11] , \U2/temp_y[10] , \U2/temp_y[9] , \U2/temp_y[8] ,
         \U2/temp_y[7] , \U2/temp_y[6] , \U2/temp_y[5] , \U2/temp_y[4] ,
         \U2/temp_y[3] , \U2/temp_y[2] , \U2/temp_y[1] , \U2/temp_y[0] ,
         \U2/temp_x[11] , \U2/temp_x[10] , \U2/temp_x[9] , \U2/temp_x[8] ,
         \U2/temp_x[7] , \U2/temp_x[6] , \U2/temp_x[5] , \U2/temp_x[4] ,
         \U2/temp_x[3] , \U2/temp_x[2] , \U2/temp_x[1] , \U2/temp_x[0] ,
         \U3/Ytt[9] , \U3/Ytt[8] , \U3/Ytt[7] , \U3/Ytt[6] , \U3/Ytt[5] ,
         \U3/Ytt[4] , \U3/Ytt[3] , \U3/Ytt[2] , \U3/Ytt[1] , \U3/Ytt[0] ,
         \U3/Xtt[9] , \U3/Xtt[8] , \U3/Xtt[7] , \U3/Xtt[6] , \U3/Xtt[5] ,
         \U3/Xtt[4] , \U3/Xtt[3] , \U3/Xtt[2] , \U3/Xtt[1] , \U3/Xtt[0] ,
         \U3/temp11[12] , \U3/temp11[1] , \U3/temp11[0] , \U3/temp12[12] ,
         \U3/temp12[1] , \U3/temp12[0] , \U3/temp10t[0] , \U3/temp10t[1] ,
         \U3/temp10t[2] , \U3/temp10t[3] , \U3/temp10t[4] , \U3/temp10t[5] ,
         \U3/temp10t[6] , \U3/temp10t[7] , \U3/temp10t[8] , \U3/temp10t[9] ,
         \U3/temp9t[0] , \U3/temp9t[1] , \U3/temp9t[2] , \U3/temp9t[3] ,
         \U3/temp9t[4] , \U3/temp9t[5] , \U3/temp9t[6] , \U3/temp9t[7] ,
         \U3/temp9t[8] , \U3/temp9t[9] , \U3/temp10[12] , \U3/temp10[11] ,
         \U3/temp9[12] , \U3/temp9[11] , \U4/Yt[11] , \U4/Yt[9] , \U4/Yt[8] ,
         \U4/Yt[7] , \U4/Yt[6] , \U4/Yt[5] , \U4/Yt[4] , \U4/Yt[3] ,
         \U4/Yt[2] , \U4/Yt[1] , \U4/Yt[0] , \U4/Xt[11] , \U4/Xt[9] ,
         \U4/Xt[8] , \U4/Xt[7] , \U4/Xt[6] , \U4/Xt[5] , \U4/Xt[4] ,
         \U4/Xt[3] , \U4/Xt[2] , \U4/Xt[1] , \U4/Xt[0] , \U4/temp7t[0] ,
         \U4/temp7t[1] , \U4/temp7t[2] , \U4/temp5t[0] , \U4/temp5t[1] ,
         \U4/temp5t[2] , \U4/temp7[11] , \U4/temp7[10] , \U4/temp7[0] ,
         \U4/temp5[11] , \U4/temp5[10] , \U4/temp5[9] , \U4/temp5[8] ,
         \U4/temp5[7] , \U4/temp5[6] , \U4/temp5[5] , \U4/temp5[4] ,
         \U4/temp5[3] , \U4/temp5[2] , \U4/temp5[1] , \U4/temp5[0] ,
         \U4/temp1[9] , \U4/temp1[7] , \U4/temp1[6] , \U4/temp1[5] ,
         \U4/temp1[4] , \U4/temp1[3] , \U4/temp1[2] , \U4/temp1[1] ,
         \U4/temp1[0] , \U4/temp2[9] , \U4/temp2[7] , \U4/temp2[6] ,
         \U4/temp2[5] , \U4/temp2[4] , \U4/temp2[3] , \U4/temp2[2] ,
         \U4/temp2[1] , \U4/temp2[0] , \U5/Yt[11] , \U5/Yt[9] , \U5/Yt[8] ,
         \U5/Yt[7] , \U5/Yt[6] , \U5/Yt[5] , \U5/Yt[4] , \U5/Yt[3] ,
         \U5/Yt[2] , \U5/Yt[1] , \U5/Yt[0] , \U5/Xt[11] , \U5/Xt[9] ,
         \U5/Xt[8] , \U5/Xt[7] , \U5/Xt[6] , \U5/Xt[5] , \U5/Xt[4] ,
         \U5/Xt[3] , \U5/Xt[2] , \U5/Xt[1] , \U5/Xt[0] , \U5/temp7t[0] ,
         \U5/temp7t[1] , \U5/temp7t[2] , \U5/temp5t[0] , \U5/temp5t[1] ,
         \U5/temp5t[2] , \U5/temp7[11] , \U5/temp7[10] , \U5/temp7[9] ,
         \U5/temp7[8] , \U5/temp7[7] , \U5/temp7[6] , \U5/temp7[5] ,
         \U5/temp7[4] , \U5/temp7[3] , \U5/temp7[2] , \U5/temp7[1] ,
         \U5/temp7[0] , \U5/temp5[11] , \U5/temp5[10] , \U5/temp5[0] ,
         \U5/temp1[9] , \U5/temp1[7] , \U5/temp1[6] , \U5/temp1[5] ,
         \U5/temp1[4] , \U5/temp1[3] , \U5/temp1[2] , \U5/temp1[1] ,
         \U5/temp1[0] , \U5/temp2[9] , \U5/temp2[7] , \U5/temp2[6] ,
         \U5/temp2[5] , \U5/temp2[4] , \U5/temp2[3] , \U5/temp2[2] ,
         \U5/temp2[1] , \U5/temp2[0] , \U6/Xt[9] , \U6/Xt[8] , \U6/Xt[7] ,
         \U6/Xt[6] , \U6/Xt[5] , \U6/Xt[4] , \U6/Xt[3] , \U6/Xt[2] ,
         \U6/Xt[1] , \U6/Xt[0] , \U6/temp6[10] , \U6/temp6[5] , \U6/temp6[4] ,
         \U6/temp6[3] , \U6/temp6[2] , \U6/temp6[1] , \U6/temp6[0] ,
         \U6/temp5[10] , \U6/temp5[5] , \U6/temp5[4] , \U6/temp5[3] ,
         \U6/temp5[2] , \U6/temp5[1] , \U6/temp5[0] , \U6/temp4t[0] ,
         \U6/temp4t[1] , \U6/temp4t[2] , \U6/temp4t[3] , \U6/temp3t[0] ,
         \U6/temp3t[1] , \U6/temp3t[2] , \U6/temp3t[3] , \U6/temp4[0] ,
         \U6/temp3[10] , \U6/temp3[9] , \U6/temp3[8] , \U6/temp3[7] ,
         \U6/temp3[6] , \U6/temp3[5] , \U6/temp3[4] , \U6/temp3[3] ,
         \U6/temp3[2] , \U6/temp3[1] , \U6/temp3[0] , \U4/U5/temp[0] ,
         \U4/U5/temp[1] , \U4/U5/temp[2] , \U4/U5/temp[3] , \U4/U5/temp[4] ,
         \U4/U5/temp[5] , \U4/U5/temp[6] , \U4/U5/temp[7] , \U4/U5/temp[11] ,
         \U4/U6/temp[0] , \U4/U6/temp[1] , \U4/U6/temp[2] , \U4/U6/temp[3] ,
         \U4/U6/temp[4] , \U4/U6/temp[5] , \U4/U6/temp[6] , \U4/U6/temp[7] ,
         \U4/U6/temp[11] , \U5/U5/temp[0] , \U5/U5/temp[1] , \U5/U5/temp[2] ,
         \U5/U5/temp[3] , \U5/U5/temp[4] , \U5/U5/temp[5] , \U5/U5/temp[6] ,
         \U5/U5/temp[7] , \U5/U5/temp[11] , \U5/U6/temp[0] , \U5/U6/temp[1] ,
         \U5/U6/temp[2] , \U5/U6/temp[3] , \U5/U6/temp[4] , \U5/U6/temp[5] ,
         \U5/U6/temp[6] , \U5/U6/temp[7] , \U5/U6/temp[11] , \intadd_25/CI ,
         \intadd_25/SUM[10] , \intadd_25/SUM[9] , \intadd_25/SUM[8] ,
         \intadd_25/SUM[7] , \intadd_25/SUM[6] , \intadd_25/SUM[5] ,
         \intadd_25/SUM[4] , \intadd_25/SUM[3] , \intadd_25/SUM[2] ,
         \intadd_25/SUM[1] , \intadd_25/SUM[0] , \intadd_25/n20 ,
         \intadd_25/n19 , \intadd_25/n18 , \intadd_25/n17 , \intadd_25/n16 ,
         \intadd_25/n15 , \intadd_25/n14 , \intadd_25/n13 , \intadd_25/n12 ,
         \intadd_25/n8 , \intadd_25/n7 , \intadd_25/n6 , \intadd_25/n5 ,
         \intadd_25/n4 , \intadd_25/n3 , \intadd_25/n2 , \intadd_26/CI ,
         \intadd_26/SUM[10] , \intadd_26/SUM[9] , \intadd_26/SUM[8] ,
         \intadd_26/SUM[7] , \intadd_26/SUM[6] , \intadd_26/SUM[5] ,
         \intadd_26/SUM[4] , \intadd_26/SUM[3] , \intadd_26/SUM[2] ,
         \intadd_26/SUM[1] , \intadd_26/SUM[0] , \intadd_26/n20 ,
         \intadd_26/n19 , \intadd_26/n18 , \intadd_26/n17 , \intadd_26/n16 ,
         \intadd_26/n15 , \intadd_26/n14 , \intadd_26/n13 , \intadd_26/n12 ,
         \intadd_26/n8 , \intadd_26/n7 , \intadd_26/n6 , \intadd_26/n5 ,
         \intadd_26/n4 , \intadd_26/n3 , \intadd_26/n2 , \intadd_29/CI ,
         \intadd_29/n11 , \intadd_29/n10 , \intadd_29/n9 , \intadd_29/n8 ,
         \intadd_29/n7 , \intadd_29/n6 , \intadd_29/n5 , \intadd_29/n4 ,
         \intadd_29/n3 , \intadd_29/n2 , \intadd_29/n1 , \intadd_30/CI ,
         \intadd_30/n11 , \intadd_30/n10 , \intadd_30/n9 , \intadd_30/n8 ,
         \intadd_30/n7 , \intadd_30/n6 , \intadd_30/n5 , \intadd_30/n4 ,
         \intadd_30/n3 , \intadd_30/n2 , \intadd_30/n1 , \intadd_31/SUM[9] ,
         \intadd_31/SUM[8] , \intadd_31/SUM[7] , \intadd_31/SUM[6] ,
         \intadd_31/SUM[5] , \intadd_31/SUM[4] , \intadd_31/SUM[3] ,
         \intadd_31/SUM[2] , \intadd_31/SUM[1] , \intadd_31/SUM[0] ,
         \intadd_31/n10 , \intadd_31/n9 , \intadd_31/n8 , \intadd_31/n7 ,
         \intadd_31/n6 , \intadd_31/n5 , \intadd_31/n4 , \intadd_31/n3 ,
         \intadd_31/n2 , \intadd_31/n1 , \intadd_32/SUM[9] ,
         \intadd_32/SUM[8] , \intadd_32/SUM[7] , \intadd_32/SUM[6] ,
         \intadd_32/SUM[5] , \intadd_32/SUM[4] , \intadd_32/SUM[3] ,
         \intadd_32/SUM[2] , \intadd_32/SUM[1] , \intadd_32/SUM[0] ,
         \intadd_32/n10 , \intadd_32/n9 , \intadd_32/n8 , \intadd_32/n7 ,
         \intadd_32/n6 , \intadd_32/n5 , \intadd_32/n4 , \intadd_32/n3 ,
         \intadd_32/n2 , \intadd_32/n1 , \intadd_34/CI , \intadd_34/n10 ,
         \intadd_34/n9 , \intadd_34/n8 , \intadd_34/n7 , \intadd_34/n6 ,
         \intadd_34/n5 , \intadd_34/n4 , \intadd_34/n3 , \intadd_34/n2 ,
         \intadd_34/n1 , \intadd_36/CI , \intadd_36/SUM[9] ,
         \intadd_36/SUM[8] , \intadd_36/SUM[7] , \intadd_36/SUM[6] ,
         \intadd_36/SUM[5] , \intadd_36/SUM[4] , \intadd_36/SUM[3] ,
         \intadd_36/SUM[2] , \intadd_36/SUM[1] , \intadd_36/SUM[0] ,
         \intadd_36/n10 , \intadd_36/n9 , \intadd_36/n8 , \intadd_36/n7 ,
         \intadd_36/n6 , \intadd_36/n5 , \intadd_36/n4 , \intadd_36/n3 ,
         \intadd_36/n2 , \intadd_36/n1 , \intadd_37/A[6] , \intadd_37/B[8] ,
         \intadd_37/B[7] , \intadd_37/B[6] , \intadd_37/B[5] ,
         \intadd_37/B[4] , \intadd_37/B[3] , \intadd_37/B[2] ,
         \intadd_37/B[1] , \intadd_37/B[0] , \intadd_37/CI , \intadd_37/n9 ,
         \intadd_37/n8 , \intadd_37/n7 , \intadd_37/n6 , \intadd_37/n5 ,
         \intadd_37/n4 , \intadd_37/n3 , \intadd_37/n2 , \intadd_37/n1 ,
         \intadd_40/CI , \intadd_40/SUM[8] , \intadd_40/SUM[7] ,
         \intadd_40/SUM[6] , \intadd_40/SUM[5] , \intadd_40/SUM[4] ,
         \intadd_40/SUM[3] , \intadd_40/SUM[2] , \intadd_40/SUM[1] ,
         \intadd_40/SUM[0] , \intadd_40/n9 , \intadd_40/n8 , \intadd_40/n7 ,
         \intadd_40/n6 , \intadd_40/n5 , \intadd_40/n4 , \intadd_40/n3 ,
         \intadd_40/n2 , \intadd_40/n1 , \intadd_41/A[8] , \intadd_41/A[7] ,
         \intadd_41/A[6] , \intadd_41/A[5] , \intadd_41/A[4] ,
         \intadd_41/A[3] , \intadd_41/A[2] , \intadd_41/A[1] ,
         \intadd_41/A[0] , \intadd_41/B[6] , \intadd_41/B[0] ,
         \intadd_41/SUM[8] , \intadd_41/SUM[7] , \intadd_41/SUM[6] ,
         \intadd_41/SUM[5] , \intadd_41/SUM[4] , \intadd_41/SUM[3] ,
         \intadd_41/SUM[2] , \intadd_41/SUM[1] , \intadd_41/SUM[0] ,
         \intadd_41/n9 , \intadd_41/n8 , \intadd_41/n7 , \intadd_41/n6 ,
         \intadd_41/n5 , \intadd_41/n4 , \intadd_41/n3 , \intadd_41/n2 ,
         \intadd_41/n1 , \intadd_49/CI , \intadd_49/n7 , \intadd_49/n6 ,
         \intadd_49/n5 , \intadd_49/n4 , \intadd_49/n3 , \intadd_49/n2 ,
         \intadd_49/n1 , \intadd_51/B[0] , \intadd_51/n3 , \intadd_51/n2 ,
         \intadd_51/n1 , \intadd_52/B[0] , \intadd_52/n3 , \intadd_52/n2 ,
         \intadd_52/n1 , \intadd_28/n1 , \intadd_33/A[6] , \intadd_33/A[5] ,
         \intadd_33/A[4] , \intadd_33/A[3] , \intadd_33/A[2] ,
         \intadd_33/A[1] , \intadd_33/A[0] , \intadd_33/SUM[9] ,
         \intadd_33/SUM[8] , \intadd_33/SUM[7] , \intadd_33/SUM[6] ,
         \intadd_33/SUM[5] , \intadd_33/SUM[4] , \intadd_33/SUM[3] ,
         \intadd_33/SUM[2] , \intadd_33/SUM[1] , \intadd_33/SUM[0] ,
         \intadd_33/n10 , \intadd_33/n9 , \intadd_33/n8 , \intadd_33/n7 ,
         \intadd_33/n6 , \intadd_33/n5 , \intadd_33/n4 , \intadd_33/n3 ,
         \intadd_33/n2 , \intadd_33/n1 , \intadd_35/A[2] , \intadd_35/A[1] ,
         \intadd_35/A[0] , \intadd_35/B[5] , \intadd_35/B[4] ,
         \intadd_35/B[3] , \intadd_35/B[2] , \intadd_35/B[1] ,
         \intadd_35/B[0] , \intadd_35/CI , \intadd_35/SUM[9] ,
         \intadd_35/SUM[8] , \intadd_35/SUM[7] , \intadd_35/SUM[6] ,
         \intadd_35/SUM[5] , \intadd_35/SUM[4] , \intadd_35/SUM[3] ,
         \intadd_35/SUM[2] , \intadd_35/SUM[1] , \intadd_35/SUM[0] ,
         \intadd_35/n10 , \intadd_35/n9 , \intadd_35/n8 , \intadd_35/n7 ,
         \intadd_35/n6 , \intadd_35/n5 , \intadd_35/n4 , \intadd_35/n3 ,
         \intadd_35/n2 , \intadd_35/n1 , \intadd_38/A[6] , \intadd_38/A[5] ,
         \intadd_38/A[4] , \intadd_38/A[3] , \intadd_38/A[2] ,
         \intadd_38/A[1] , \intadd_38/A[0] , \intadd_38/B[7] ,
         \intadd_38/B[6] , \intadd_38/B[5] , \intadd_38/B[4] ,
         \intadd_38/B[3] , \intadd_38/B[2] , \intadd_38/B[1] ,
         \intadd_38/B[0] , \intadd_38/CI , \intadd_38/SUM[8] ,
         \intadd_38/SUM[7] , \intadd_38/SUM[6] , \intadd_38/SUM[5] ,
         \intadd_38/SUM[4] , \intadd_38/SUM[3] , \intadd_38/SUM[2] ,
         \intadd_38/SUM[1] , \intadd_38/SUM[0] , \intadd_38/n9 ,
         \intadd_38/n8 , \intadd_38/n7 , \intadd_38/n6 , \intadd_38/n5 ,
         \intadd_38/n4 , \intadd_38/n3 , \intadd_38/n2 , \intadd_38/n1 ,
         \intadd_39/A[1] , \intadd_39/A[0] , \intadd_39/B[8] ,
         \intadd_39/B[7] , \intadd_39/B[6] , \intadd_39/B[5] ,
         \intadd_39/B[4] , \intadd_39/B[3] , \intadd_39/B[2] ,
         \intadd_39/B[1] , \intadd_39/CI , \intadd_39/n9 , \intadd_39/n8 ,
         \intadd_39/n7 , \intadd_39/n6 , \intadd_39/n5 , \intadd_39/n4 ,
         \intadd_39/n3 , \intadd_39/n2 , \intadd_39/n1 , \intadd_42/A[2] ,
         \intadd_42/A[1] , \intadd_42/A[0] , \intadd_42/B[6] ,
         \intadd_42/B[0] , \intadd_42/n9 , \intadd_42/n8 , \intadd_42/n7 ,
         \intadd_42/n6 , \intadd_42/n5 , \intadd_42/n4 , \intadd_42/n3 ,
         \intadd_42/n2 , \intadd_42/n1 , \intadd_43/A[7] , \intadd_43/A[1] ,
         \intadd_43/B[5] , \intadd_43/B[3] , \intadd_43/B[1] ,
         \intadd_43/B[0] , \intadd_43/CI , \intadd_43/n9 , \intadd_43/n8 ,
         \intadd_43/n7 , \intadd_43/n6 , \intadd_43/n5 , \intadd_43/n4 ,
         \intadd_43/n3 , \intadd_43/n2 , \intadd_43/n1 , \intadd_44/A[7] ,
         \intadd_44/A[1] , \intadd_44/B[3] , \intadd_44/B[1] ,
         \intadd_44/B[0] , \intadd_44/CI , \intadd_44/n9 , \intadd_44/n8 ,
         \intadd_44/n7 , \intadd_44/n6 , \intadd_44/n5 , \intadd_44/n4 ,
         \intadd_44/n3 , \intadd_44/n2 , \intadd_44/n1 , \intadd_45/A[8] ,
         \intadd_45/B[0] , \intadd_45/CI , \intadd_45/SUM[2] ,
         \intadd_45/SUM[1] , \intadd_45/SUM[0] , \intadd_45/n9 ,
         \intadd_45/n8 , \intadd_45/n7 , \intadd_45/n6 , \intadd_45/n5 ,
         \intadd_45/n4 , \intadd_45/n3 , \intadd_45/n2 , \intadd_45/n1 ,
         \intadd_46/CI , \intadd_46/n8 , \intadd_46/n7 , \intadd_46/n6 ,
         \intadd_46/n5 , \intadd_46/n4 , \intadd_46/n3 , \intadd_46/n2 ,
         \intadd_46/n1 , \intadd_47/CI , \intadd_47/n8 , \intadd_47/n7 ,
         \intadd_47/n6 , \intadd_47/n5 , \intadd_47/n4 , \intadd_47/n3 ,
         \intadd_47/n2 , \intadd_47/n1 , \intadd_48/CI , \intadd_48/n8 ,
         \intadd_48/n7 , \intadd_48/n6 , \intadd_48/n5 , \intadd_48/n4 ,
         \intadd_48/n3 , \intadd_48/n2 , \intadd_48/n1 , \intadd_50/CI ,
         \intadd_50/n7 , \intadd_50/n6 , \intadd_50/n5 , \intadd_50/n4 ,
         \intadd_50/n3 , \intadd_50/n2 , \intadd_50/n1 , n561, n562, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, n623,
         n625, n626, n627, n628, n630, n631, n632, n633, n635, n636, n637,
         n638, n639, n640, n643, n646, n649, n650, n651, n652, n654, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n702, n703, n704, n705,
         n706, n707, n708, n710, n711, n712, n714, n715, n716, n718, n719,
         n720, n721, n723, n724, n725, n726, n727, n728, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n743, n744, n745,
         n746, n747, n748, n749, n751, n752, n754, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n973, n974, n975,
         n976, n977, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1001, n1002, n1003, n1005, n1006, n1007, n1008, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1066, n1067, n1069, n1071, n1072, n1074, n1077, n1079,
         n1080, n1081, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1110, n1111, n1112,
         n1113, n1114, n1115, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1302, n1303, n1305, n1306, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1354, n1355, n1357, n1358, n1360, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1405, n1406, n1407,
         n1408, n1409, n1411, n1412, n1413, n1414, n1415, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1458, n1459, n1460, n1461, n1463, n1464, n1467, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1486, n1487, n1488, n1489, n1490, n1493,
         n1494, n1495, n1496, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1515,
         n1516, n1517, n1518, n1519, n1520, n1633, n1635, n1638, n1639, n1640,
         n1641, n1642, n1643, n1645, n1646, n1647, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1660, n1661, n1662, n1664,
         n1666, n1668, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1713, n1714, n1715, n1716, n1717, n1719,
         n1721, n1722, n1725, n1726, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1780, n1781, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1793,
         n1795, n1796, n1797, n1798, n1799, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1856, n1859, n1860, n1862,
         n1865, n1867, n1868, n1870, n1871, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1884, n1885, n1886, n1887, n1888,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1959, n1961, n1962, n1964, n1965,
         n1966, n1968, n1969, n1972, n1973, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2004, n2005, n2006, n2007, n2008, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n1883, n1637, n1644, n1648, n1724, n1790, n1741, n1728, n2020,
         n1659, n1770, n1855, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844;
  wire   [9:0] temp1;
  wire   [9:0] temp2;
  wire   [9:0] temp3;
  wire   [9:0] temp4;
  wire   [9:0] temp5;
  wire   [9:0] temp6;
  wire   [9:0] temp7;
  wire   [9:0] temp8;
  wire   [9:0] temp1t;
  wire   [9:0] temp2t;
  wire   [9:0] temp3t;
  wire   [9:0] temp4t;
  wire   [12:0] s0;
  wire   [12:0] s1;
  wire   [12:0] s2;
  wire   [12:0] s3;
  wire   [11:0] result1;
  wire   [11:0] result2;
  wire   [11:0] result3;
  wire   [11:0] result4;
  wire   [11:0] result5;
  wire   [11:0] result6;
  wire   [11:0] result7;
  wire   [11:0] result8;
  wire   [12:0] s4;
  wire   [12:0] s5;
  assign D2[12] = D2[10];
  assign D2[11] = D2[10];
  assign D3[11] = D3[12];
  assign D5[11] = D5[12];
  assign D6[12] = D6[10];
  assign D6[11] = D6[10];

  DFFHQX4 \U11/temp_reg[0]  ( .D(temp4[0]), .CK(clk), .Q(\temp5t[0] ) );
  DFFHQX4 \U11/temp_reg[1]  ( .D(temp5[1]), .CK(clk), .Q(\U5/temp1[0] ) );
  DFFHQX4 \U12/temp_reg[0]  ( .D(temp3[0]), .CK(clk), .Q(\temp6t[0] ) );
  DFFHQX4 \U13/temp_reg[0]  ( .D(temp2[0]), .CK(clk), .Q(\temp7t[0] ) );
  DFFHQX4 \U14/temp_reg[0]  ( .D(temp1[0]), .CK(clk), .Q(\temp8t[0] ) );
  DFFHQX1 \U16/temp_reg[0]  ( .D(s4[0]), .CK(clk), .Q(D1[0]) );
  DFFHQX1 \U16/temp_reg[1]  ( .D(s4[1]), .CK(clk), .Q(D1[1]) );
  DFFHQX1 \U16/temp_reg[2]  ( .D(s4[2]), .CK(clk), .Q(D1[2]) );
  DFFHQX1 \U16/temp_reg[3]  ( .D(s4[3]), .CK(clk), .Q(D1[3]) );
  DFFHQX1 \U16/temp_reg[4]  ( .D(s4[4]), .CK(clk), .Q(D1[4]) );
  DFFHQX1 \U16/temp_reg[5]  ( .D(s4[5]), .CK(clk), .Q(D1[5]) );
  DFFHQX1 \U16/temp_reg[6]  ( .D(s4[6]), .CK(clk), .Q(D1[6]) );
  DFFHQX1 \U16/temp_reg[7]  ( .D(s4[7]), .CK(clk), .Q(D1[7]) );
  DFFHQX1 \U16/temp_reg[8]  ( .D(s4[8]), .CK(clk), .Q(D1[8]) );
  DFFHQX1 \U16/temp_reg[9]  ( .D(s4[9]), .CK(clk), .Q(D1[9]) );
  DFFHQX1 \U16/temp_reg[10]  ( .D(s4[10]), .CK(clk), .Q(D1[10]) );
  DFFHQX1 \U16/temp_reg[11]  ( .D(s4[11]), .CK(clk), .Q(D1[11]) );
  DFFHQX1 \U16/temp_reg[12]  ( .D(n853), .CK(clk), .Q(D1[12]) );
  DFFHQX1 \U18/temp_reg[0]  ( .D(\s6[0] ), .CK(clk), .Q(D3[0]) );
  DFFHQX1 \U18/temp_reg[1]  ( .D(n914), .CK(clk), .Q(D3[1]) );
  DFFHQX1 \U18/temp_reg[2]  ( .D(n908), .CK(clk), .Q(D3[2]) );
  DFFHQX1 \U18/temp_reg[3]  ( .D(n894), .CK(clk), .Q(D3[3]) );
  DFFHQX1 \U18/temp_reg[4]  ( .D(n893), .CK(clk), .Q(D3[4]) );
  DFFHQX1 \U18/temp_reg[5]  ( .D(n886), .CK(clk), .Q(D3[5]) );
  DFFHQX1 \U18/temp_reg[6]  ( .D(n870), .CK(clk), .Q(D3[6]) );
  DFFHQX1 \U18/temp_reg[7]  ( .D(n869), .CK(clk), .Q(D3[7]) );
  DFFHQX1 \U18/temp_reg[8]  ( .D(n865), .CK(clk), .Q(D3[8]) );
  DFFHQX1 \U18/temp_reg[9]  ( .D(n858), .CK(clk), .Q(D3[9]) );
  DFFHQX1 \U18/temp_reg[10]  ( .D(n857), .CK(clk), .Q(D3[10]) );
  DFFHQX1 \U20/temp_reg[0]  ( .D(\s7[0] ), .CK(clk), .Q(D5[0]) );
  DFFHQX1 \U20/temp_reg[1]  ( .D(n917), .CK(clk), .Q(D5[1]) );
  DFFHQX1 \U20/temp_reg[2]  ( .D(n909), .CK(clk), .Q(D5[2]) );
  DFFHQX1 \U20/temp_reg[3]  ( .D(n899), .CK(clk), .Q(D5[3]) );
  DFFHQX1 \U20/temp_reg[4]  ( .D(n898), .CK(clk), .Q(D5[4]) );
  DFFHQX1 \U20/temp_reg[5]  ( .D(n887), .CK(clk), .Q(D5[5]) );
  DFFHQX1 \U20/temp_reg[6]  ( .D(n875), .CK(clk), .Q(D5[6]) );
  DFFHQX1 \U20/temp_reg[7]  ( .D(n874), .CK(clk), .Q(D5[7]) );
  DFFHQX1 \U20/temp_reg[8]  ( .D(n866), .CK(clk), .Q(D5[8]) );
  DFFHQX1 \U20/temp_reg[9]  ( .D(n861), .CK(clk), .Q(D5[9]) );
  DFFHQX1 \U20/temp_reg[10]  ( .D(n860), .CK(clk), .Q(D5[10]) );
  DFFHQX1 \U22/temp_reg[0]  ( .D(s5[0]), .CK(clk), .Q(D7[0]) );
  DFFHQX1 \U22/temp_reg[1]  ( .D(s5[1]), .CK(clk), .Q(D7[1]) );
  DFFHQX1 \U22/temp_reg[2]  ( .D(s5[2]), .CK(clk), .Q(D7[2]) );
  DFFHQX1 \U22/temp_reg[3]  ( .D(s5[3]), .CK(clk), .Q(D7[3]) );
  DFFHQX1 \U22/temp_reg[4]  ( .D(s5[4]), .CK(clk), .Q(D7[4]) );
  DFFHQX1 \U22/temp_reg[5]  ( .D(s5[5]), .CK(clk), .Q(D7[5]) );
  DFFHQX1 \U22/temp_reg[6]  ( .D(s5[6]), .CK(clk), .Q(D7[6]) );
  DFFHQX1 \U22/temp_reg[7]  ( .D(s5[7]), .CK(clk), .Q(D7[7]) );
  DFFHQX1 \U22/temp_reg[8]  ( .D(s5[8]), .CK(clk), .Q(D7[8]) );
  DFFHQX1 \U22/temp_reg[9]  ( .D(s5[9]), .CK(clk), .Q(D7[9]) );
  DFFHQX1 \U22/temp_reg[10]  ( .D(s5[10]), .CK(clk), .Q(D7[10]) );
  DFFHQX1 \U22/temp_reg[11]  ( .D(s5[11]), .CK(clk), .Q(D7[11]) );
  DFFHQX1 \U22/temp_reg[12]  ( .D(n855), .CK(clk), .Q(D7[12]) );
  DFFHQX1 \U19/temp_reg[0]  ( .D(s0[0]), .CK(clk), .Q(D4[0]) );
  DFFHQX1 \U19/temp_reg[1]  ( .D(s0[1]), .CK(clk), .Q(D4[1]) );
  DFFHQX1 \U19/temp_reg[2]  ( .D(s0[2]), .CK(clk), .Q(D4[2]) );
  DFFHQX1 \U19/temp_reg[3]  ( .D(s0[3]), .CK(clk), .Q(D4[3]) );
  DFFHQX1 \U19/temp_reg[4]  ( .D(s0[4]), .CK(clk), .Q(D4[4]) );
  DFFHQX1 \U19/temp_reg[5]  ( .D(s0[5]), .CK(clk), .Q(D4[5]) );
  DFFHQX1 \U19/temp_reg[6]  ( .D(s0[6]), .CK(clk), .Q(D4[6]) );
  DFFHQX1 \U19/temp_reg[7]  ( .D(s0[7]), .CK(clk), .Q(D4[7]) );
  DFFHQX1 \U19/temp_reg[8]  ( .D(s0[8]), .CK(clk), .Q(D4[8]) );
  DFFHQX1 \U19/temp_reg[9]  ( .D(s0[9]), .CK(clk), .Q(D4[9]) );
  DFFHQX1 \U19/temp_reg[10]  ( .D(s0[10]), .CK(clk), .Q(D4[10]) );
  DFFHQX1 \U19/temp_reg[11]  ( .D(s0[11]), .CK(clk), .Q(D4[11]) );
  DFFHQX1 \U19/temp_reg[12]  ( .D(s0[12]), .CK(clk), .Q(D4[12]) );
  DFFHQX1 \U15/temp_reg[0]  ( .D(s1[0]), .CK(clk), .Q(D0[0]) );
  DFFHQX1 \U15/temp_reg[1]  ( .D(s1[1]), .CK(clk), .Q(D0[1]) );
  DFFHQX1 \U15/temp_reg[2]  ( .D(s1[2]), .CK(clk), .Q(D0[2]) );
  DFFHQX1 \U15/temp_reg[3]  ( .D(s1[3]), .CK(clk), .Q(D0[3]) );
  DFFHQX1 \U15/temp_reg[4]  ( .D(s1[4]), .CK(clk), .Q(D0[4]) );
  DFFHQX1 \U15/temp_reg[5]  ( .D(s1[5]), .CK(clk), .Q(D0[5]) );
  DFFHQX1 \U15/temp_reg[6]  ( .D(s1[6]), .CK(clk), .Q(D0[6]) );
  DFFHQX1 \U15/temp_reg[7]  ( .D(s1[7]), .CK(clk), .Q(D0[7]) );
  DFFHQX1 \U15/temp_reg[8]  ( .D(s1[8]), .CK(clk), .Q(D0[8]) );
  DFFHQX1 \U15/temp_reg[9]  ( .D(s1[9]), .CK(clk), .Q(D0[9]) );
  DFFHQX1 \U15/temp_reg[10]  ( .D(s1[10]), .CK(clk), .Q(D0[10]) );
  DFFHQX1 \U15/temp_reg[11]  ( .D(s1[11]), .CK(clk), .Q(D0[11]) );
  DFFHQX1 \U15/temp_reg[12]  ( .D(s1[12]), .CK(clk), .Q(D0[12]) );
  DFFHQX1 \U21/temp_reg[0]  ( .D(s2[0]), .CK(clk), .Q(D6[0]) );
  DFFHQX1 \U21/temp_reg[1]  ( .D(s2[1]), .CK(clk), .Q(D6[1]) );
  DFFHQX1 \U21/temp_reg[2]  ( .D(s2[2]), .CK(clk), .Q(D6[2]) );
  DFFHQX1 \U21/temp_reg[3]  ( .D(s2[3]), .CK(clk), .Q(D6[3]) );
  DFFHQX1 \U21/temp_reg[4]  ( .D(s2[4]), .CK(clk), .Q(D6[4]) );
  DFFHQX1 \U21/temp_reg[5]  ( .D(s2[5]), .CK(clk), .Q(D6[5]) );
  DFFHQX1 \U21/temp_reg[6]  ( .D(s2[6]), .CK(clk), .Q(D6[6]) );
  DFFHQX1 \U21/temp_reg[7]  ( .D(s2[7]), .CK(clk), .Q(D6[7]) );
  DFFHQX1 \U21/temp_reg[8]  ( .D(s2[8]), .CK(clk), .Q(D6[8]) );
  DFFHQX1 \U21/temp_reg[9]  ( .D(s2[9]), .CK(clk), .Q(D6[9]) );
  DFFHQX1 \U17/temp_reg[0]  ( .D(s3[0]), .CK(clk), .Q(D2[0]) );
  DFFHQX1 \U17/temp_reg[1]  ( .D(s3[1]), .CK(clk), .Q(D2[1]) );
  DFFHQX1 \U17/temp_reg[2]  ( .D(s3[2]), .CK(clk), .Q(D2[2]) );
  DFFHQX1 \U17/temp_reg[3]  ( .D(s3[3]), .CK(clk), .Q(D2[3]) );
  DFFHQX1 \U17/temp_reg[4]  ( .D(s3[4]), .CK(clk), .Q(D2[4]) );
  DFFHQX1 \U17/temp_reg[5]  ( .D(s3[5]), .CK(clk), .Q(D2[5]) );
  DFFHQX1 \U17/temp_reg[6]  ( .D(s3[6]), .CK(clk), .Q(D2[6]) );
  DFFHQX1 \U17/temp_reg[7]  ( .D(s3[7]), .CK(clk), .Q(D2[7]) );
  DFFHQX1 \U17/temp_reg[8]  ( .D(s3[8]), .CK(clk), .Q(D2[8]) );
  DFFHQX1 \U17/temp_reg[9]  ( .D(s3[9]), .CK(clk), .Q(D2[9]) );
  DFFHQX1 \U18/temp_reg[12]  ( .D(\intadd_31/n1 ), .CK(clk), .Q(D3[12]) );
  DFFHQX1 \U20/temp_reg[12]  ( .D(\intadd_32/n1 ), .CK(clk), .Q(D5[12]) );
  DFFHQX1 \U21/temp_reg[10]  ( .D(s2[12]), .CK(clk), .Q(D6[10]) );
  DFFHQX1 \U17/temp_reg[10]  ( .D(s3[12]), .CK(clk), .Q(D2[10]) );
  DFFHQX1 \U1/U22/temp_reg[0]  ( .D(\U1/Xtt[0] ), .CK(clk), .Q(s0[0]) );
  DFFHQX1 \U1/U22/temp_reg[1]  ( .D(\U1/Xtt[1] ), .CK(clk), .Q(s0[1]) );
  DFFHQX1 \U1/U22/temp_reg[2]  ( .D(\U1/Xtt[2] ), .CK(clk), .Q(s0[2]) );
  DFFHQX1 \U1/U22/temp_reg[3]  ( .D(\U1/Xtt[3] ), .CK(clk), .Q(s0[3]) );
  DFFHQX1 \U1/U22/temp_reg[4]  ( .D(\U1/Xtt[4] ), .CK(clk), .Q(s0[4]) );
  DFFHQX1 \U1/U22/temp_reg[5]  ( .D(\U1/Xtt[5] ), .CK(clk), .Q(s0[5]) );
  DFFHQX1 \U1/U22/temp_reg[6]  ( .D(\U1/Xtt[6] ), .CK(clk), .Q(s0[6]) );
  DFFHQX1 \U1/U22/temp_reg[7]  ( .D(\U1/Xtt[7] ), .CK(clk), .Q(s0[7]) );
  DFFHQX1 \U1/U22/temp_reg[8]  ( .D(\U1/Xtt[8] ), .CK(clk), .Q(s0[8]) );
  DFFHQX1 \U1/U22/temp_reg[9]  ( .D(\U1/Xtt[9] ), .CK(clk), .Q(s0[9]) );
  DFFHQX1 \U1/U22/temp_reg[10]  ( .D(\U1/Xtt[10] ), .CK(clk), .Q(s0[10]) );
  DFFHQX1 \U1/U22/temp_reg[11]  ( .D(\U1/Xtt[11] ), .CK(clk), .Q(s0[11]) );
  DFFHQX1 \U1/U22/temp_reg[12]  ( .D(\U1/result5[13] ), .CK(clk), .Q(s0[12])
         );
  DFFHQX1 \U1/U23/temp_reg[0]  ( .D(\U1/Ytt[0] ), .CK(clk), .Q(s1[0]) );
  DFFHQX1 \U1/U23/temp_reg[1]  ( .D(\U1/Ytt[1] ), .CK(clk), .Q(s1[1]) );
  DFFHQX1 \U1/U23/temp_reg[2]  ( .D(\U1/Ytt[2] ), .CK(clk), .Q(s1[2]) );
  DFFHQX1 \U1/U23/temp_reg[3]  ( .D(\U1/Ytt[3] ), .CK(clk), .Q(s1[3]) );
  DFFHQX1 \U1/U23/temp_reg[4]  ( .D(\U1/Ytt[4] ), .CK(clk), .Q(s1[4]) );
  DFFHQX1 \U1/U23/temp_reg[5]  ( .D(\U1/Ytt[5] ), .CK(clk), .Q(s1[5]) );
  DFFHQX1 \U1/U23/temp_reg[6]  ( .D(\U1/Ytt[6] ), .CK(clk), .Q(s1[6]) );
  DFFHQX1 \U1/U23/temp_reg[7]  ( .D(\U1/Ytt[7] ), .CK(clk), .Q(s1[7]) );
  DFFHQX1 \U1/U23/temp_reg[8]  ( .D(\U1/Ytt[8] ), .CK(clk), .Q(s1[8]) );
  DFFHQX1 \U1/U23/temp_reg[9]  ( .D(\U1/Ytt[9] ), .CK(clk), .Q(s1[9]) );
  DFFHQX1 \U1/U23/temp_reg[10]  ( .D(\U1/Ytt[10] ), .CK(clk), .Q(s1[10]) );
  DFFHQX1 \U1/U23/temp_reg[11]  ( .D(\U1/Ytt[11] ), .CK(clk), .Q(s1[11]) );
  DFFHQX1 \U1/U23/temp_reg[12]  ( .D(\U1/result6[13] ), .CK(clk), .Q(s1[12])
         );
  DFFHQX1 \U2/U22/temp_reg[0]  ( .D(\U2/Xtt[0] ), .CK(clk), .Q(s2[0]) );
  DFFHQX1 \U2/U22/temp_reg[1]  ( .D(\U2/Xtt[1] ), .CK(clk), .Q(s2[1]) );
  DFFHQX1 \U2/U22/temp_reg[2]  ( .D(\U2/Xtt[2] ), .CK(clk), .Q(s2[2]) );
  DFFHQX1 \U2/U22/temp_reg[3]  ( .D(\U2/Xtt[3] ), .CK(clk), .Q(s2[3]) );
  DFFHQX1 \U2/U22/temp_reg[4]  ( .D(\U2/Xtt[4] ), .CK(clk), .Q(s2[4]) );
  DFFHQX1 \U2/U22/temp_reg[5]  ( .D(\U2/Xtt[5] ), .CK(clk), .Q(s2[5]) );
  DFFHQX1 \U2/U22/temp_reg[6]  ( .D(\U2/Xtt[6] ), .CK(clk), .Q(s2[6]) );
  DFFHQX1 \U2/U22/temp_reg[7]  ( .D(\U2/Xtt[7] ), .CK(clk), .Q(s2[7]) );
  DFFHQX1 \U2/U22/temp_reg[8]  ( .D(\U2/Xtt[8] ), .CK(clk), .Q(s2[8]) );
  DFFHQX1 \U2/U22/temp_reg[9]  ( .D(\U2/Xtt[9] ), .CK(clk), .Q(s2[9]) );
  DFFHQX1 \U2/U22/temp_reg[12]  ( .D(\U2/Xtt[10] ), .CK(clk), .Q(s2[12]) );
  DFFHQX1 \U2/U23/temp_reg[0]  ( .D(\U2/Ytt[0] ), .CK(clk), .Q(s3[0]) );
  DFFHQX1 \U2/U23/temp_reg[1]  ( .D(\U2/Ytt[1] ), .CK(clk), .Q(s3[1]) );
  DFFHQX1 \U2/U23/temp_reg[2]  ( .D(\U2/Ytt[2] ), .CK(clk), .Q(s3[2]) );
  DFFHQX1 \U2/U23/temp_reg[3]  ( .D(\U2/Ytt[3] ), .CK(clk), .Q(s3[3]) );
  DFFHQX1 \U2/U23/temp_reg[4]  ( .D(\U2/Ytt[4] ), .CK(clk), .Q(s3[4]) );
  DFFHQX1 \U2/U23/temp_reg[5]  ( .D(\U2/Ytt[5] ), .CK(clk), .Q(s3[5]) );
  DFFHQX1 \U2/U23/temp_reg[6]  ( .D(\U2/Ytt[6] ), .CK(clk), .Q(s3[6]) );
  DFFHQX1 \U2/U23/temp_reg[7]  ( .D(\U2/Ytt[7] ), .CK(clk), .Q(s3[7]) );
  DFFHQX1 \U2/U23/temp_reg[8]  ( .D(\U2/Ytt[8] ), .CK(clk), .Q(s3[8]) );
  DFFHQX1 \U2/U23/temp_reg[9]  ( .D(\U2/Ytt[9] ), .CK(clk), .Q(s3[9]) );
  DFFHQX1 \U2/U23/temp_reg[12]  ( .D(\U2/Ytt[10] ), .CK(clk), .Q(s3[12]) );
  DFFHQX1 \U3/U22/temp_reg[11]  ( .D(n2842), .CK(clk), .Q(result1[11]) );
  DFFHQX1 \U3/U23/temp_reg[11]  ( .D(\intadd_28/n1 ), .CK(clk), .Q(result2[11]) );
  DFFHQX1 \U5/U13/temp_reg[9]  ( .D(\U5/Xt[9] ), .CK(clk), .Q(result5[9]) );
  DFFHQX1 \U5/U14/temp_reg[9]  ( .D(\U5/Yt[9] ), .CK(clk), .Q(result6[9]) );
  DFFHQX1 \U6/U9/temp_reg[11]  ( .D(n884), .CK(clk), .Q(result7[11]) );
  DFFHQX1 \U6/U10/temp_reg[11]  ( .D(\intadd_36/n1 ), .CK(clk), .Q(result8[11]) );
  DFFHQX1 \U3/U22/temp_reg[9]  ( .D(\U3/Xtt[9] ), .CK(clk), .Q(result1[9]) );
  DFFHQX1 \U3/U22/temp_reg[10]  ( .D(n2843), .CK(clk), .Q(result1[10]) );
  DFFHQX1 \U3/U23/temp_reg[9]  ( .D(\U3/Ytt[9] ), .CK(clk), .Q(result2[9]) );
  DFFHQX1 \U3/U23/temp_reg[10]  ( .D(n2844), .CK(clk), .Q(result2[10]) );
  DFFHQX1 \U4/U13/temp_reg[9]  ( .D(\U4/Xt[9] ), .CK(clk), .Q(result3[9]) );
  DFFHQX1 \U5/U14/temp_reg[11]  ( .D(\U5/Yt[11] ), .CK(clk), .Q(result6[11])
         );
  DFFHQX1 \U6/U9/temp_reg[8]  ( .D(\U6/Xt[8] ), .CK(clk), .Q(result7[8]) );
  DFFHQX1 \U6/U9/temp_reg[9]  ( .D(\U6/Xt[9] ), .CK(clk), .Q(result7[9]) );
  DFFHQX1 \U6/U10/temp_reg[8]  ( .D(n880), .CK(clk), .Q(result8[8]) );
  DFFHQX1 \U6/U10/temp_reg[9]  ( .D(n879), .CK(clk), .Q(result8[9]) );
  DFFHQX1 \U4/U13/temp_reg[11]  ( .D(\U4/Xt[11] ), .CK(clk), .Q(result3[11])
         );
  DFFHQX1 \U4/U14/temp_reg[11]  ( .D(\U4/Yt[11] ), .CK(clk), .Q(result4[11])
         );
  DFFHQX1 \U5/U13/temp_reg[6]  ( .D(\U5/Xt[6] ), .CK(clk), .Q(result5[6]) );
  DFFHQX1 \U5/U13/temp_reg[7]  ( .D(\U5/Xt[7] ), .CK(clk), .Q(result5[7]) );
  DFFHQX1 \U5/U13/temp_reg[8]  ( .D(\U5/Xt[8] ), .CK(clk), .Q(result5[8]) );
  DFFHQX1 \U5/U14/temp_reg[6]  ( .D(\U5/Yt[6] ), .CK(clk), .Q(result6[6]) );
  DFFHQX1 \U5/U14/temp_reg[7]  ( .D(\U5/Yt[7] ), .CK(clk), .Q(result6[7]) );
  DFFHQX1 \U5/U14/temp_reg[8]  ( .D(\U5/Yt[8] ), .CK(clk), .Q(result6[8]) );
  DFFHQX1 \U6/U7/temp_reg[10]  ( .D(\U6/temp3[10] ), .CK(clk), .Q(
        \U6/temp5[10] ) );
  DFFHQX1 \U3/U22/temp_reg[6]  ( .D(\U3/Xtt[6] ), .CK(clk), .Q(result1[6]) );
  DFFHQX1 \U3/U22/temp_reg[7]  ( .D(\U3/Xtt[7] ), .CK(clk), .Q(result1[7]) );
  DFFHQX1 \U3/U22/temp_reg[8]  ( .D(\U3/Xtt[8] ), .CK(clk), .Q(result1[8]) );
  DFFHQX1 \U3/U23/temp_reg[6]  ( .D(\U3/Ytt[6] ), .CK(clk), .Q(result2[6]) );
  DFFHQX1 \U3/U23/temp_reg[7]  ( .D(\U3/Ytt[7] ), .CK(clk), .Q(result2[7]) );
  DFFHQX1 \U3/U23/temp_reg[8]  ( .D(\U3/Ytt[8] ), .CK(clk), .Q(result2[8]) );
  DFFHQX1 \U4/U13/temp_reg[5]  ( .D(\U4/Xt[5] ), .CK(clk), .Q(result3[5]) );
  DFFHQX1 \U4/U13/temp_reg[6]  ( .D(\U4/Xt[6] ), .CK(clk), .Q(result3[6]) );
  DFFHQX1 \U4/U13/temp_reg[7]  ( .D(\U4/Xt[7] ), .CK(clk), .Q(result3[7]) );
  DFFHQX1 \U4/U14/temp_reg[5]  ( .D(\U4/Yt[5] ), .CK(clk), .Q(result4[5]) );
  DFFHQX1 \U4/U14/temp_reg[6]  ( .D(\U4/Yt[6] ), .CK(clk), .Q(result4[6]) );
  DFFHQX1 \U4/U14/temp_reg[7]  ( .D(\U4/Yt[7] ), .CK(clk), .Q(result4[7]) );
  DFFHQX1 \U4/U14/temp_reg[8]  ( .D(\U4/Yt[8] ), .CK(clk), .Q(result4[8]) );
  DFFHQX1 \U6/U9/temp_reg[5]  ( .D(\U6/Xt[5] ), .CK(clk), .Q(result7[5]) );
  DFFHQX1 \U6/U9/temp_reg[6]  ( .D(\U6/Xt[6] ), .CK(clk), .Q(result7[6]) );
  DFFHQX1 \U6/U9/temp_reg[7]  ( .D(\U6/Xt[7] ), .CK(clk), .Q(result7[7]) );
  DFFHQX1 \U6/U10/temp_reg[5]  ( .D(n883), .CK(clk), .Q(result8[5]) );
  DFFHQX1 \U6/U10/temp_reg[6]  ( .D(n882), .CK(clk), .Q(result8[6]) );
  DFFHQX1 \U6/U10/temp_reg[7]  ( .D(n881), .CK(clk), .Q(result8[7]) );
  DFFHQX1 \U6/U7/temp_reg[9]  ( .D(\U6/temp3[9] ), .CK(clk), .Q(\U6/temp5[5] )
         );
  DFFHQX1 \U6/U8/temp_reg[9]  ( .D(n839), .CK(clk), .Q(\U6/temp6[5] ) );
  DFFHQX1 \U2/U21/temp_reg[9]  ( .D(\U2/temp_y[9] ), .CK(clk), .Q(
        \U2/result2[8] ) );
  DFFHQX1 \U5/U13/temp_reg[3]  ( .D(\U5/Xt[3] ), .CK(clk), .Q(result5[3]) );
  DFFHQX1 \U5/U13/temp_reg[4]  ( .D(\U5/Xt[4] ), .CK(clk), .Q(result5[4]) );
  DFFHQX1 \U5/U13/temp_reg[5]  ( .D(\U5/Xt[5] ), .CK(clk), .Q(result5[5]) );
  DFFHQX1 \U5/U14/temp_reg[3]  ( .D(\U5/Yt[3] ), .CK(clk), .Q(result6[3]) );
  DFFHQX1 \U5/U14/temp_reg[4]  ( .D(\U5/Yt[4] ), .CK(clk), .Q(result6[4]) );
  DFFHQX1 \U5/U14/temp_reg[5]  ( .D(\U5/Yt[5] ), .CK(clk), .Q(result6[5]) );
  DFFHQX1 \U6/U8/temp_reg[2]  ( .D(n846), .CK(clk), .Q(\U6/temp4t[2] ) );
  DFFHQX1 \U6/U8/temp_reg[3]  ( .D(n845), .CK(clk), .Q(\U6/temp4t[3] ) );
  DFFHQX1 \U3/U22/temp_reg[2]  ( .D(\U3/Xtt[2] ), .CK(clk), .Q(result1[2]) );
  DFFHQX1 \U3/U22/temp_reg[3]  ( .D(\U3/Xtt[3] ), .CK(clk), .Q(result1[3]) );
  DFFHQX1 \U3/U22/temp_reg[4]  ( .D(\U3/Xtt[4] ), .CK(clk), .Q(result1[4]) );
  DFFHQX1 \U3/U22/temp_reg[5]  ( .D(\U3/Xtt[5] ), .CK(clk), .Q(result1[5]) );
  DFFHQX1 \U3/U23/temp_reg[2]  ( .D(\U3/Ytt[2] ), .CK(clk), .Q(result2[2]) );
  DFFHQX1 \U3/U23/temp_reg[3]  ( .D(\U3/Ytt[3] ), .CK(clk), .Q(result2[3]) );
  DFFHQX1 \U3/U23/temp_reg[4]  ( .D(\U3/Ytt[4] ), .CK(clk), .Q(result2[4]) );
  DFFHQX1 \U3/U23/temp_reg[5]  ( .D(\U3/Ytt[5] ), .CK(clk), .Q(result2[5]) );
  DFFHQX1 \U6/U7/temp_reg[1]  ( .D(\U6/temp3[1] ), .CK(clk), .Q(\U6/temp3t[1] ) );
  DFFHQX1 \U6/U7/temp_reg[2]  ( .D(\U6/temp3[2] ), .CK(clk), .Q(\U6/temp3t[2] ) );
  DFFHQX1 \U6/U7/temp_reg[3]  ( .D(\U6/temp3[3] ), .CK(clk), .Q(\U6/temp3t[3] ) );
  DFFHQX1 \U4/U13/temp_reg[2]  ( .D(\U4/Xt[2] ), .CK(clk), .Q(result3[2]) );
  DFFHQX1 \U4/U13/temp_reg[3]  ( .D(\U4/Xt[3] ), .CK(clk), .Q(result3[3]) );
  DFFHQX1 \U4/U13/temp_reg[4]  ( .D(\U4/Xt[4] ), .CK(clk), .Q(result3[4]) );
  DFFHQX1 \U4/U14/temp_reg[2]  ( .D(\U4/Yt[2] ), .CK(clk), .Q(result4[2]) );
  DFFHQX1 \U4/U14/temp_reg[3]  ( .D(\U4/Yt[3] ), .CK(clk), .Q(result4[3]) );
  DFFHQX1 \U4/U14/temp_reg[4]  ( .D(\U4/Yt[4] ), .CK(clk), .Q(result4[4]) );
  DFFHQX1 \U6/U9/temp_reg[2]  ( .D(\U6/Xt[2] ), .CK(clk), .Q(result7[2]) );
  DFFHQX1 \U6/U9/temp_reg[3]  ( .D(\U6/Xt[3] ), .CK(clk), .Q(result7[3]) );
  DFFHQX1 \U6/U9/temp_reg[4]  ( .D(\U6/Xt[4] ), .CK(clk), .Q(result7[4]) );
  DFFHQX1 \U6/U10/temp_reg[2]  ( .D(n904), .CK(clk), .Q(result8[2]) );
  DFFHQX1 \U6/U10/temp_reg[3]  ( .D(n903), .CK(clk), .Q(result8[3]) );
  DFFHQX1 \U6/U10/temp_reg[4]  ( .D(n890), .CK(clk), .Q(result8[4]) );
  DFFHQX1 \U6/U7/temp_reg[6]  ( .D(\U6/temp3[6] ), .CK(clk), .Q(\U6/temp5[2] )
         );
  DFFHQX1 \U6/U7/temp_reg[7]  ( .D(\U6/temp3[7] ), .CK(clk), .Q(\U6/temp5[3] )
         );
  DFFHQX1 \U6/U7/temp_reg[8]  ( .D(\U6/temp3[8] ), .CK(clk), .Q(\U6/temp5[4] )
         );
  DFFHQX1 \U2/U21/temp_reg[8]  ( .D(\U2/temp_y[8] ), .CK(clk), .Q(
        \U2/result2[7] ) );
  DFFHQX1 \U6/U8/temp_reg[6]  ( .D(n842), .CK(clk), .Q(\U6/temp6[2] ) );
  DFFHQX1 \U6/U8/temp_reg[7]  ( .D(n841), .CK(clk), .Q(\U6/temp6[3] ) );
  DFFHQX1 \U6/U8/temp_reg[8]  ( .D(n840), .CK(clk), .Q(\U6/temp6[4] ) );
  DFFHQX1 \U6/U7/temp_reg[0]  ( .D(\U6/temp3[0] ), .CK(clk), .Q(\U6/temp3t[0] ) );
  DFFHQX1 \U2/U20/temp_reg[9]  ( .D(\U2/temp_x[9] ), .CK(clk), .Q(
        \U2/result1[8] ) );
  DFFHQX1 \U5/U13/temp_reg[1]  ( .D(\U5/Xt[1] ), .CK(clk), .Q(result5[1]) );
  DFFHQX1 \U5/U13/temp_reg[2]  ( .D(\U5/Xt[2] ), .CK(clk), .Q(result5[2]) );
  DFFHQX1 \U5/U14/temp_reg[1]  ( .D(\U5/Yt[1] ), .CK(clk), .Q(result6[1]) );
  DFFHQX1 \U5/U14/temp_reg[2]  ( .D(\U5/Yt[2] ), .CK(clk), .Q(result6[2]) );
  DFFHQX1 \U6/U8/temp_reg[1]  ( .D(n847), .CK(clk), .Q(\U6/temp4t[1] ) );
  DFFHQX1 \U6/U8/temp_reg[0]  ( .D(\U6/temp4[0] ), .CK(clk), .Q(\U6/temp4t[0] ) );
  DFFHQX1 \U3/U22/temp_reg[1]  ( .D(\U3/Xtt[1] ), .CK(clk), .Q(result1[1]) );
  DFFHQX1 \U3/U23/temp_reg[1]  ( .D(\U3/Ytt[1] ), .CK(clk), .Q(result2[1]) );
  DFFHQX1 \U4/U13/temp_reg[1]  ( .D(\U4/Xt[1] ), .CK(clk), .Q(result3[1]) );
  DFFHQX1 \U4/U14/temp_reg[1]  ( .D(\U4/Yt[1] ), .CK(clk), .Q(result4[1]) );
  DFFHQX1 \U6/U9/temp_reg[1]  ( .D(\U6/Xt[1] ), .CK(clk), .Q(result7[1]) );
  DFFHQX1 \U6/U10/temp_reg[1]  ( .D(n905), .CK(clk), .Q(result8[1]) );
  DFFHQX1 \U4/U13/temp_reg[0]  ( .D(\U4/Xt[0] ), .CK(clk), .Q(result3[0]) );
  DFFHQX1 \U4/U14/temp_reg[0]  ( .D(\U4/Yt[0] ), .CK(clk), .Q(result4[0]) );
  DFFHQX1 \U3/U22/temp_reg[0]  ( .D(\U3/Xtt[0] ), .CK(clk), .Q(result1[0]) );
  DFFHQX1 \U3/U23/temp_reg[0]  ( .D(\U3/Ytt[0] ), .CK(clk), .Q(result2[0]) );
  DFFHQX1 \U6/U8/temp_reg[4]  ( .D(n844), .CK(clk), .Q(\U6/temp6[0] ) );
  DFFHQX1 \U6/U9/temp_reg[0]  ( .D(\U6/Xt[0] ), .CK(clk), .Q(result7[0]) );
  DFFHQX1 \U6/U10/temp_reg[0]  ( .D(n920), .CK(clk), .Q(result8[0]) );
  DFFHQX1 \U6/U7/temp_reg[4]  ( .D(\U6/temp3[4] ), .CK(clk), .Q(\U6/temp5[0] )
         );
  DFFHQX1 \U6/U8/temp_reg[5]  ( .D(n843), .CK(clk), .Q(\U6/temp6[1] ) );
  DFFHQX1 \U6/U7/temp_reg[5]  ( .D(\U6/temp3[5] ), .CK(clk), .Q(\U6/temp5[1] )
         );
  DFFHQX1 \U2/U20/temp_reg[8]  ( .D(\U2/temp_x[8] ), .CK(clk), .Q(
        \U2/result1[7] ) );
  DFFHQX1 \U2/U20/temp_reg[7]  ( .D(\U2/temp_x[7] ), .CK(clk), .Q(
        \U2/result1[6] ) );
  DFFHQX1 \U2/U21/temp_reg[7]  ( .D(\U2/temp_y[7] ), .CK(clk), .Q(
        \U2/result2[6] ) );
  DFFHQX1 \U5/U13/temp_reg[0]  ( .D(\U5/Xt[0] ), .CK(clk), .Q(result5[0]) );
  DFFHQX1 \U5/U14/temp_reg[0]  ( .D(\U5/Yt[0] ), .CK(clk), .Q(result6[0]) );
  DFFHQX1 \U2/U21/temp_reg[6]  ( .D(\U2/temp_y[6] ), .CK(clk), .Q(
        \U2/result2[5] ) );
  DFFHQX1 \U12/temp_reg[7]  ( .D(temp6[7]), .CK(clk), .Q(\U4/temp1[6] ) );
  DFFHQX1 \U13/temp_reg[8]  ( .D(temp7[8]), .CK(clk), .Q(\U4/temp2[7] ) );
  DFFHQX1 \U2/U20/temp_reg[5]  ( .D(\U2/temp_x[5] ), .CK(clk), .Q(
        \U2/result1[4] ) );
  DFFHQX1 \U2/U21/temp_reg[5]  ( .D(\U2/temp_y[5] ), .CK(clk), .Q(
        \U2/result2[4] ) );
  DFFHQX1 \U1/U20/temp_reg[7]  ( .D(\U1/temp_xxx[7] ), .CK(clk), .Q(
        \U1/temp_xxxt[7] ) );
  DFFHQX1 \U1/U21/temp_reg[7]  ( .D(\U1/temp_yyy[7] ), .CK(clk), .Q(
        \U1/temp_yyyt[7] ) );
  DFFHQX1 \U3/U20/temp_reg[7]  ( .D(n684), .CK(clk), .Q(\U3/temp9t[7] ) );
  DFFHQX1 \U3/U20/temp_reg[8]  ( .D(n683), .CK(clk), .Q(\U3/temp9t[8] ) );
  DFFHQX1 \U3/U20/temp_reg[9]  ( .D(n682), .CK(clk), .Q(\U3/temp9t[9] ) );
  DFFHQX1 \U2/U20/temp_reg[6]  ( .D(\U2/temp_x[6] ), .CK(clk), .Q(
        \U2/result1[5] ) );
  DFFHQX1 \U7/temp_reg[8]  ( .D(temp1[8]), .CK(clk), .Q(temp1t[8]) );
  DFFHQX1 \U8/temp_reg[8]  ( .D(temp2[8]), .CK(clk), .Q(temp2t[8]) );
  DFFHQX1 \U10/temp_reg[7]  ( .D(temp4[7]), .CK(clk), .Q(temp4t[7]) );
  DFFHQX1 \U4/U11/temp_reg[10]  ( .D(\U4/temp5[10] ), .CK(clk), .Q(
        \U4/U5/temp[7] ) );
  DFFHQX1 \U4/U12/temp_reg[10]  ( .D(\U4/temp7[10] ), .CK(clk), .Q(
        \U4/U6/temp[7] ) );
  DFFHQX1 \U5/U11/temp_reg[10]  ( .D(\U5/temp5[10] ), .CK(clk), .Q(
        \U5/U5/temp[7] ) );
  DFFHQX1 \U5/U12/temp_reg[10]  ( .D(\U5/temp7[10] ), .CK(clk), .Q(
        \U5/U6/temp[7] ) );
  DFFHQX1 \U10/temp_reg[9]  ( .D(temp4[9]), .CK(clk), .Q(temp4t[9]) );
  DFFHQX1 \U8/temp_reg[9]  ( .D(temp2[9]), .CK(clk), .Q(temp2t[9]) );
  DFFHQX1 \U14/temp_reg[8]  ( .D(temp8[8]), .CK(clk), .Q(\U5/temp2[7] ) );
  DFFHQX1 \U13/temp_reg[4]  ( .D(temp7[4]), .CK(clk), .Q(\U4/temp2[3] ) );
  DFFHQX1 \U13/temp_reg[5]  ( .D(temp7[5]), .CK(clk), .Q(\U4/temp2[4] ) );
  DFFHQX1 \U12/temp_reg[6]  ( .D(temp6[6]), .CK(clk), .Q(\U4/temp1[5] ) );
  DFFHQX1 \U12/temp_reg[4]  ( .D(temp6[4]), .CK(clk), .Q(\U4/temp1[3] ) );
  DFFHQX1 \U12/temp_reg[5]  ( .D(temp6[5]), .CK(clk), .Q(\U4/temp1[4] ) );
  DFFHQX1 \U13/temp_reg[7]  ( .D(temp7[7]), .CK(clk), .Q(\U4/temp2[6] ) );
  DFFHQX1 \U13/temp_reg[6]  ( .D(temp7[6]), .CK(clk), .Q(\U4/temp2[5] ) );
  DFFHQX1 \U1/U20/temp_reg[4]  ( .D(\U1/temp_xxx[4] ), .CK(clk), .Q(
        \U1/temp_xxxt[4] ) );
  DFFHQX1 \U1/U21/temp_reg[4]  ( .D(\U1/temp_yyy[4] ), .CK(clk), .Q(
        \U1/temp_yyyt[4] ) );
  DFFHQX1 \U1/U20/temp_reg[5]  ( .D(\U1/temp_xxx[5] ), .CK(clk), .Q(
        \U1/temp_xxxt[5] ) );
  DFFHQX1 \U1/U20/temp_reg[6]  ( .D(\U1/temp_xxx[6] ), .CK(clk), .Q(
        \U1/temp_xxxt[6] ) );
  DFFHQX1 \U1/U21/temp_reg[5]  ( .D(\U1/temp_yyy[5] ), .CK(clk), .Q(
        \U1/temp_yyyt[5] ) );
  DFFHQX1 \U1/U21/temp_reg[6]  ( .D(\U1/temp_yyy[6] ), .CK(clk), .Q(
        \U1/temp_yyyt[6] ) );
  DFFHQX1 \U3/U20/temp_reg[4]  ( .D(n698), .CK(clk), .Q(\U3/temp9t[4] ) );
  DFFHQX1 \U3/U20/temp_reg[5]  ( .D(n697), .CK(clk), .Q(\U3/temp9t[5] ) );
  DFFHQX1 \U3/U20/temp_reg[6]  ( .D(n693), .CK(clk), .Q(\U3/temp9t[6] ) );
  DFFHQX1 \U2/U20/temp_reg[4]  ( .D(\U2/temp_x[4] ), .CK(clk), .Q(
        \U2/result1[3] ) );
  DFFHQX1 \U2/U21/temp_reg[4]  ( .D(\U2/temp_y[4] ), .CK(clk), .Q(
        \U2/result2[3] ) );
  DFFHQX1 \U7/temp_reg[6]  ( .D(temp1[6]), .CK(clk), .Q(temp1t[6]) );
  DFFHQX1 \U8/temp_reg[4]  ( .D(temp2[4]), .CK(clk), .Q(temp2t[4]) );
  DFFHQX1 \U8/temp_reg[6]  ( .D(temp2[6]), .CK(clk), .Q(temp2t[6]) );
  DFFHQX1 \U8/temp_reg[7]  ( .D(temp2[7]), .CK(clk), .Q(temp2t[7]) );
  DFFHQX1 \U9/temp_reg[5]  ( .D(temp3[5]), .CK(clk), .Q(temp3t[5]) );
  DFFHQX1 \U9/temp_reg[6]  ( .D(temp3[6]), .CK(clk), .Q(temp3t[6]) );
  DFFHQX1 \U9/temp_reg[7]  ( .D(temp3[7]), .CK(clk), .Q(temp3t[7]) );
  DFFHQX1 \U10/temp_reg[5]  ( .D(temp4[5]), .CK(clk), .Q(temp4t[5]) );
  DFFHQX1 \U4/U11/temp_reg[6]  ( .D(\U4/temp5[6] ), .CK(clk), .Q(
        \U4/U5/temp[3] ) );
  DFFHQX1 \U4/U11/temp_reg[8]  ( .D(\U4/temp5[8] ), .CK(clk), .Q(
        \U4/U5/temp[5] ) );
  DFFHQX1 \U4/U12/temp_reg[6]  ( .D(n816), .CK(clk), .Q(\U4/U6/temp[3] ) );
  DFFHQX1 \U4/U12/temp_reg[8]  ( .D(n814), .CK(clk), .Q(\U4/U6/temp[5] ) );
  DFFHQX1 \U5/U11/temp_reg[6]  ( .D(n792), .CK(clk), .Q(\U5/U5/temp[3] ) );
  DFFHQX1 \U5/U11/temp_reg[8]  ( .D(n790), .CK(clk), .Q(\U5/U5/temp[5] ) );
  DFFHQX1 \U5/U12/temp_reg[6]  ( .D(\U5/temp7[6] ), .CK(clk), .Q(
        \U5/U6/temp[3] ) );
  DFFHQX1 \U5/U12/temp_reg[8]  ( .D(\U5/temp7[8] ), .CK(clk), .Q(
        \U5/U6/temp[5] ) );
  DFFHQX1 \U13/temp_reg[1]  ( .D(temp7[1]), .CK(clk), .Q(\U4/temp2[0] ) );
  DFFHQX1 \U11/temp_reg[8]  ( .D(temp5[8]), .CK(clk), .Q(\U5/temp1[7] ) );
  DFFHQX1 \U13/temp_reg[2]  ( .D(temp7[2]), .CK(clk), .Q(\U4/temp2[1] ) );
  DFFHQX1 \U13/temp_reg[3]  ( .D(temp7[3]), .CK(clk), .Q(\U4/temp2[2] ) );
  DFFHQX1 \U12/temp_reg[2]  ( .D(temp6[2]), .CK(clk), .Q(\U4/temp1[1] ) );
  DFFHQX1 \U14/temp_reg[6]  ( .D(temp8[6]), .CK(clk), .Q(\U5/temp2[5] ) );
  DFFHQX1 \U12/temp_reg[3]  ( .D(temp6[3]), .CK(clk), .Q(\U4/temp1[2] ) );
  DFFHQX1 \U3/U21/temp_reg[1]  ( .D(n716), .CK(clk), .Q(\U3/temp10t[1] ) );
  DFFHQX1 \U1/U20/temp_reg[1]  ( .D(\U1/temp_xxx[1] ), .CK(clk), .Q(
        \U1/temp_xxxt[1] ) );
  DFFHQX1 \U1/U20/temp_reg[2]  ( .D(\U1/temp_xxx[2] ), .CK(clk), .Q(
        \U1/temp_xxxt[2] ) );
  DFFHQX1 \U1/U20/temp_reg[3]  ( .D(\U1/temp_xxx[3] ), .CK(clk), .Q(
        \U1/temp_xxxt[3] ) );
  DFFHQX1 \U1/U21/temp_reg[1]  ( .D(\U1/temp_yyy[1] ), .CK(clk), .Q(
        \U1/temp_yyyt[1] ) );
  DFFHQX1 \U1/U21/temp_reg[2]  ( .D(\U1/temp_yyy[2] ), .CK(clk), .Q(
        \U1/temp_yyyt[2] ) );
  DFFHQX1 \U1/U21/temp_reg[3]  ( .D(\U1/temp_yyy[3] ), .CK(clk), .Q(
        \U1/temp_yyyt[3] ) );
  DFFHQX1 \U3/U20/temp_reg[1]  ( .D(n710), .CK(clk), .Q(\U3/temp9t[1] ) );
  DFFHQX1 \U4/U11/temp_reg[2]  ( .D(\U4/temp5[2] ), .CK(clk), .Q(
        \U4/temp5t[2] ) );
  DFFHQX1 \U4/U12/temp_reg[1]  ( .D(n821), .CK(clk), .Q(\U4/temp7t[1] ) );
  DFFHQX1 \U4/U12/temp_reg[2]  ( .D(n820), .CK(clk), .Q(\U4/temp7t[2] ) );
  DFFHQX1 \U5/U11/temp_reg[2]  ( .D(n797), .CK(clk), .Q(\U5/temp5t[2] ) );
  DFFHQX1 \U5/U12/temp_reg[2]  ( .D(\U5/temp7[2] ), .CK(clk), .Q(
        \U5/temp7t[2] ) );
  DFFHQX1 \U3/U20/temp_reg[2]  ( .D(n706), .CK(clk), .Q(\U3/temp9t[2] ) );
  DFFHQX1 \U3/U20/temp_reg[3]  ( .D(n702), .CK(clk), .Q(\U3/temp9t[3] ) );
  DFFHQX1 \U3/U20/temp_reg[12]  ( .D(\U3/temp9[12] ), .CK(clk), .Q(
        \U3/temp12[12] ) );
  DFFHQX1 \U3/U21/temp_reg[0]  ( .D(n2051), .CK(clk), .Q(\U3/temp10t[0] ) );
  DFFHQX1 \U4/U11/temp_reg[1]  ( .D(\U4/temp5[1] ), .CK(clk), .Q(
        \U4/temp5t[1] ) );
  DFFHQX1 \U5/U11/temp_reg[1]  ( .D(n798), .CK(clk), .Q(\U5/temp5t[1] ) );
  DFFHQX1 \U3/U20/temp_reg[10]  ( .D(n681), .CK(clk), .Q(\U3/temp12[0] ) );
  DFFHQX1 \U9/temp_reg[3]  ( .D(temp3[3]), .CK(clk), .Q(temp3t[3]) );
  DFFHQX1 \U10/temp_reg[3]  ( .D(temp4[3]), .CK(clk), .Q(temp4t[3]) );
  DFFHQX1 \U4/U11/temp_reg[4]  ( .D(\U4/temp5[4] ), .CK(clk), .Q(
        \U4/U5/temp[1] ) );
  DFFHQX1 \U4/U12/temp_reg[4]  ( .D(n818), .CK(clk), .Q(\U4/U6/temp[1] ) );
  DFFHQX1 \U5/U11/temp_reg[4]  ( .D(n795), .CK(clk), .Q(\U5/U5/temp[1] ) );
  DFFHQX1 \U5/U12/temp_reg[4]  ( .D(\U5/temp7[4] ), .CK(clk), .Q(
        \U5/U6/temp[1] ) );
  DFFHQX1 \U5/U11/temp_reg[0]  ( .D(\U5/temp5[0] ), .CK(clk), .Q(
        \U5/temp5t[0] ) );
  DFFHQX1 \U11/temp_reg[6]  ( .D(temp5[6]), .CK(clk), .Q(\U5/temp1[5] ) );
  DFFHQX1 \U14/temp_reg[7]  ( .D(temp8[7]), .CK(clk), .Q(\U5/temp2[6] ) );
  DFFHQX1 \U14/temp_reg[4]  ( .D(temp8[4]), .CK(clk), .Q(\U5/temp2[3] ) );
  DFFHQX1 \U3/U20/temp_reg[0]  ( .D(n2049), .CK(clk), .Q(\U3/temp9t[0] ) );
  DFFHQX1 \U2/U20/temp_reg[3]  ( .D(\U2/temp_x[3] ), .CK(clk), .Q(
        \U2/result1[2] ) );
  DFFHQX1 \U2/U21/temp_reg[3]  ( .D(\U2/temp_y[3] ), .CK(clk), .Q(
        \U2/result2[2] ) );
  DFFHQX1 \U1/U20/temp_reg[0]  ( .D(\U1/temp_xxx[0] ), .CK(clk), .Q(
        \U1/temp_xxxt[0] ) );
  DFFHQX1 \U1/U21/temp_reg[0]  ( .D(n649), .CK(clk), .Q(\U1/temp_yyyt[0] ) );
  DFFHQX1 \U2/U20/temp_reg[2]  ( .D(\U2/temp_x[2] ), .CK(clk), .Q(
        \U2/result1[1] ) );
  DFFHQX1 \U2/U21/temp_reg[2]  ( .D(\U2/temp_y[2] ), .CK(clk), .Q(
        \U2/result2[1] ) );
  DFFHQX1 \U2/U20/temp_reg[1]  ( .D(\U2/temp_x[1] ), .CK(clk), .Q(
        \U2/result1[0] ) );
  DFFHQX1 \U2/U21/temp_reg[1]  ( .D(\U2/temp_y[1] ), .CK(clk), .Q(
        \U2/result2[0] ) );
  DFFHQX1 \U2/U20/temp_reg[0]  ( .D(\U2/temp_x[0] ), .CK(clk), .Q(
        \U2/temp_xt[0] ) );
  DFFHQX1 \U2/U21/temp_reg[0]  ( .D(\U2/temp_y[0] ), .CK(clk), .Q(
        \U2/temp_yt[0] ) );
  DFFHQX1 \U12/temp_reg[1]  ( .D(temp6[1]), .CK(clk), .Q(\U4/temp1[0] ) );
  DFFHQX1 \U11/temp_reg[4]  ( .D(temp5[4]), .CK(clk), .Q(\U5/temp1[3] ) );
  DFFHQX4 \U1/U21/temp_reg[13]  ( .D(\U1/temp_yyy[11] ), .CK(clk), .Q(
        \U1/result6[13] ) );
  DFFHQX4 \U1/U20/temp_reg[13]  ( .D(\U1/temp_xxx[11] ), .CK(clk), .Q(
        \U1/result5[13] ) );
  AOI222X1 U572 ( .A0(x7[8]), .A1(n561), .B0(x7[8]), .B1(n1126), .C0(n561), 
        .C1(n1126), .Y(temp8[9]) );
  AOI2BB2X1 U587 ( .B0(n1141), .B1(n1140), .A0N(n1140), .A1N(n1141), .Y(
        temp8[1]) );
  AOI2BB2X1 U603 ( .B0(n1157), .B1(n1156), .A0N(n1156), .A1N(n1157), .Y(
        temp7[1]) );
  AOI222X1 U604 ( .A0(x5[8]), .A1(n589), .B0(x5[8]), .B1(n1158), .C0(n589), 
        .C1(n1158), .Y(temp6[9]) );
  AOI2BB2X1 U619 ( .B0(n1173), .B1(n1172), .A0N(n1172), .A1N(n1173), .Y(
        temp6[1]) );
  AOI2BB2X1 U635 ( .B0(n1189), .B1(n1188), .A0N(n1188), .A1N(n1189), .Y(
        temp5[1]) );
  OAI21XL U636 ( .A0(n617), .A1(n603), .B0(n1190), .Y(temp4[9]) );
  OAI21XL U662 ( .A0(x4[0]), .A1(n616), .B0(n1188), .Y(temp4[0]) );
  OAI21XL U664 ( .A0(n622), .A1(n589), .B0(n1199), .Y(temp3[9]) );
  OAI21XL U690 ( .A0(x5[0]), .A1(n602), .B0(n1172), .Y(temp3[0]) );
  OAI21XL U692 ( .A0(n627), .A1(n575), .B0(n1208), .Y(temp2[9]) );
  OAI21XL U718 ( .A0(x6[0]), .A1(n588), .B0(n1156), .Y(temp2[0]) );
  OAI21XL U720 ( .A0(n632), .A1(n561), .B0(n1217), .Y(temp1[9]) );
  OAI21XL U721 ( .A0(x7[8]), .A1(x0[8]), .B0(n1218), .Y(n1217) );
  OAI21XL U746 ( .A0(x7[0]), .A1(n574), .B0(n1140), .Y(temp1[0]) );
  OAI21XL U748 ( .A0(result8[0]), .A1(n933), .B0(n1226), .Y(\s7[0] ) );
  OAI21XL U749 ( .A0(result7[0]), .A1(n932), .B0(n1227), .Y(\s6[0] ) );
  AOI22X1 U750 ( .A0(result4[0]), .A1(result2[0]), .B0(n925), .B1(n923), .Y(
        s5[0]) );
  AOI22X1 U751 ( .A0(result3[0]), .A1(result1[0]), .B0(n924), .B1(n922), .Y(
        s4[0]) );
  AOI21X1 U754 ( .A0(n764), .A1(n1230), .B0(n2050), .Y(n1229) );
  AOI21X1 U766 ( .A0(n1240), .A1(n1230), .B0(\intadd_45/CI ), .Y(n1239) );
  NOR2X1 U771 ( .A(n812), .B(n1058), .Y(\intadd_49/CI ) );
  AOI2BB1X1 U777 ( .A0N(\U2/result2[1] ), .A1N(n1250), .B0(n1104), .Y(
        \intadd_44/CI ) );
  AOI211X1 U781 ( .A0(n1108), .A1(n1106), .B0(n1250), .C0(n1102), .Y(
        \intadd_44/B[0] ) );
  NOR2X1 U782 ( .A(n1108), .B(n1106), .Y(n1250) );
  AOI22X1 U784 ( .A0(n1104), .A1(\U2/result2[2] ), .B0(n1102), .B1(n1255), .Y(
        \intadd_44/A[1] ) );
  AOI2BB1X1 U785 ( .A0N(\U2/result1[1] ), .A1N(n1256), .B0(n1103), .Y(
        \intadd_43/CI ) );
  AOI211X1 U789 ( .A0(n1107), .A1(n1105), .B0(n1256), .C0(n1101), .Y(
        \intadd_43/B[0] ) );
  NOR2X1 U790 ( .A(n1107), .B(n1105), .Y(n1256) );
  NAND2BX1 U791 ( .AN(\U2/Xtt[10] ), .B(n1260), .Y(\intadd_43/A[7] ) );
  AOI22X1 U792 ( .A0(n1103), .A1(\U2/result1[2] ), .B0(n1101), .B1(n1261), .Y(
        \intadd_43/A[1] ) );
  NOR2X1 U798 ( .A(\temp7t[0] ), .B(n1061), .Y(\intadd_40/CI ) );
  OAI2BB2X1 U816 ( .B0(n1281), .B1(n1267), .A0N(n1267), .A1N(n1281), .Y(
        \intadd_39/A[1] ) );
  AOI22X1 U818 ( .A0(n2551), .A1(n1230), .B0(n801), .B1(n787), .Y(
        \intadd_39/A[0] ) );
  NOR2BX1 U823 ( .AN(\U6/temp5[0] ), .B(\U6/temp4t[0] ), .Y(\intadd_36/CI ) );
  NOR2BX1 U829 ( .AN(\U6/temp3t[0] ), .B(n926), .Y(\intadd_34/CI ) );
  AOI22X1 U838 ( .A0(\temp7t[0] ), .A1(\U4/temp1[2] ), .B0(n1061), .B1(n850), 
        .Y(\U6/temp4[0] ) );
  AOI2BB1X1 U840 ( .A0N(n811), .A1N(n1287), .B0(n1288), .Y(n1286) );
  AOI22X1 U842 ( .A0(\intadd_49/n1 ), .A1(n1289), .B0(n1113), .B1(n811), .Y(
        \U6/temp3[8] ) );
  AOI21X1 U844 ( .A0(n1290), .A1(n1119), .B0(n1291), .Y(\U6/temp3[10] ) );
  AOI21X1 U845 ( .A0(\U4/temp1[9] ), .A1(n1265), .B0(n811), .Y(n1291) );
  NAND2X1 U846 ( .A(\U4/temp1[7] ), .B(n1114), .Y(n1265) );
  NAND2X1 U847 ( .A(\U4/temp2[9] ), .B(n1118), .Y(n1290) );
  AOI22X1 U848 ( .A0(n2568), .A1(\U4/temp2[2] ), .B0(n1058), .B1(n812), .Y(
        \U6/temp3[0] ) );
  AOI222X1 U849 ( .A0(n803), .A1(n793), .B0(n803), .B1(\intadd_42/n1 ), .C0(
        n793), .C1(\intadd_42/n1 ), .Y(\U5/temp7[11] ) );
  OAI21XL U854 ( .A0(n803), .A1(\intadd_38/A[6] ), .B0(n1293), .Y(
        \U5/temp5[11] ) );
  OAI21XL U855 ( .A0(n793), .A1(\intadd_42/B[6] ), .B0(\intadd_38/n1 ), .Y(
        n1293) );
  NOR2X1 U862 ( .A(\U5/temp1[0] ), .B(n851), .Y(n1299) );
  MXI2X1 U871 ( .A(n1302), .B(n2137), .S0(n1309), .Y(\U5/Yt[6] ) );
  AOI2BB2X1 U872 ( .B0(n1008), .B1(n1310), .A0N(n1310), .A1N(n1008), .Y(n1309)
         );
  MXI2X1 U873 ( .A(n1302), .B(n2137), .S0(n1311), .Y(\U5/Yt[5] ) );
  AOI2BB2X1 U874 ( .B0(n1312), .B1(n1313), .A0N(n1312), .A1N(n1313), .Y(n1311)
         );
  MXI2X1 U875 ( .A(n1302), .B(n2137), .S0(n1314), .Y(\U5/Yt[4] ) );
  AOI2BB2X1 U876 ( .B0(n1315), .B1(n1316), .A0N(n1316), .A1N(n1315), .Y(n1314)
         );
  AOI22X1 U891 ( .A0(\U5/U6/temp[4] ), .A1(\U5/U6/temp[1] ), .B0(n1092), .B1(
        n1053), .Y(n1329) );
  AOI22X1 U893 ( .A0(\U5/U6/temp[11] ), .A1(\U5/U6/temp[7] ), .B0(n1010), .B1(
        n1022), .Y(n1331) );
  AOI22X1 U900 ( .A0(\U5/U6/temp[2] ), .A1(\U5/temp7t[2] ), .B0(n1074), .B1(
        n1093), .Y(n1334) );
  AOI22X1 U903 ( .A0(\U5/U6/temp[11] ), .A1(n1054), .B0(\U5/U6/temp[5] ), .B1(
        n1022), .Y(n1336) );
  AOI2BB2X1 U910 ( .B0(\U5/U6/temp[0] ), .B1(n1052), .A0N(n1052), .A1N(
        \U5/U6/temp[0] ), .Y(n1340) );
  AOI22X1 U912 ( .A0(\U5/U6/temp[5] ), .A1(n1093), .B0(\U5/U6/temp[2] ), .B1(
        n1054), .Y(n1342) );
  AOI2BB2X1 U921 ( .B0(\U5/temp7t[1] ), .B1(n1092), .A0N(n1092), .A1N(
        \U5/temp7t[1] ), .Y(n1347) );
  AOI22X1 U925 ( .A0(\U5/U6/temp[6] ), .A1(n1052), .B0(\U5/U6/temp[3] ), .B1(
        n1007), .Y(n1350) );
  AOI22X1 U927 ( .A0(\U5/U6/temp[7] ), .A1(n1053), .B0(\U5/U6/temp[4] ), .B1(
        n1010), .Y(n1351) );
  AOI2BB2X1 U944 ( .B0(n1364), .B1(n1365), .A0N(n1364), .A1N(n1365), .Y(n1363)
         );
  AOI2BB2X1 U946 ( .B0(n1367), .B1(n1368), .A0N(n1368), .A1N(n1367), .Y(n1366)
         );
  AOI22X1 U961 ( .A0(\U5/U5/temp[4] ), .A1(\U5/U5/temp[1] ), .B0(n1090), .B1(
        n1050), .Y(n1381) );
  AOI22X1 U963 ( .A0(\U5/U5/temp[11] ), .A1(\U5/U5/temp[7] ), .B0(n998), .B1(
        n1021), .Y(n1383) );
  AOI22X1 U968 ( .A0(\U5/U5/temp[2] ), .A1(\U5/temp5t[2] ), .B0(n1071), .B1(
        n1091), .Y(n1386) );
  AOI22X1 U970 ( .A0(\U5/U5/temp[11] ), .A1(n1051), .B0(\U5/U5/temp[5] ), .B1(
        n1021), .Y(n1388) );
  AOI2BB2X1 U973 ( .B0(\U5/U5/temp[0] ), .B1(n1049), .A0N(n1049), .A1N(
        \U5/U5/temp[0] ), .Y(n1392) );
  AOI22X1 U975 ( .A0(\U5/U5/temp[5] ), .A1(n1091), .B0(\U5/U5/temp[2] ), .B1(
        n1051), .Y(n1394) );
  AOI22X1 U977 ( .A0(\U5/U5/temp[11] ), .A1(n995), .B0(\U5/U5/temp[6] ), .B1(
        n1021), .Y(n1395) );
  AOI2BB2X1 U984 ( .B0(\U5/temp5t[1] ), .B1(n1090), .A0N(n1090), .A1N(
        \U5/temp5t[1] ), .Y(n1399) );
  AOI22X1 U988 ( .A0(\U5/U5/temp[6] ), .A1(n1049), .B0(\U5/U5/temp[3] ), .B1(
        n995), .Y(n1402) );
  OAI21XL U998 ( .A0(n825), .A1(\intadd_41/B[6] ), .B0(n1404), .Y(
        \U4/temp7[11] ) );
  OAI21XL U999 ( .A0(n848), .A1(\intadd_37/A[6] ), .B0(\intadd_41/n1 ), .Y(
        n1404) );
  AOI21X1 U1002 ( .A0(\intadd_50/CI ), .A1(n849), .B0(\intadd_41/B[0] ), .Y(
        n1407) );
  AOI211X1 U1003 ( .A0(n2568), .A1(n1055), .B0(\intadd_50/CI ), .C0(n849), .Y(
        \intadd_41/B[0] ) );
  NAND2X1 U1005 ( .A(n2568), .B(n1055), .Y(n1406) );
  AOI222X1 U1006 ( .A0(n848), .A1(\intadd_37/n1 ), .B0(n848), .B1(n825), .C0(
        \intadd_37/n1 ), .C1(n825), .Y(\U4/temp5[11] ) );
  AOI2BB2X1 U1026 ( .B0(n1421), .B1(n1422), .A0N(n1421), .A1N(n1422), .Y(n1420) );
  AOI2BB2X1 U1028 ( .B0(n1424), .B1(n1425), .A0N(n1425), .A1N(n1424), .Y(n1423) );
  AOI2BB2X1 U1032 ( .B0(n1430), .B1(n1431), .A0N(n1431), .A1N(n1430), .Y(n1429) );
  AOI22X1 U1043 ( .A0(\U4/U6/temp[4] ), .A1(\U4/U6/temp[1] ), .B0(n1088), .B1(
        n1047), .Y(n1438) );
  AOI22X1 U1045 ( .A0(\U4/U6/temp[11] ), .A1(\U4/U6/temp[7] ), .B0(n986), .B1(
        n1020), .Y(n1440) );
  AOI22X1 U1050 ( .A0(\U4/U6/temp[2] ), .A1(\U4/temp7t[2] ), .B0(n1069), .B1(
        n1089), .Y(n1443) );
  AOI2BB2X1 U1055 ( .B0(\U4/U6/temp[0] ), .B1(n1046), .A0N(n1046), .A1N(
        \U4/U6/temp[0] ), .Y(n1449) );
  AOI22X1 U1057 ( .A0(\U4/U6/temp[5] ), .A1(n1089), .B0(\U4/U6/temp[2] ), .B1(
        n1048), .Y(n1451) );
  AOI22X1 U1059 ( .A0(\U4/U6/temp[11] ), .A1(n983), .B0(\U4/U6/temp[6] ), .B1(
        n1020), .Y(n1452) );
  AOI2BB2X1 U1066 ( .B0(\U4/temp7t[1] ), .B1(n1088), .A0N(n1088), .A1N(
        \U4/temp7t[1] ), .Y(n1456) );
  AOI22X1 U1070 ( .A0(\U4/U6/temp[6] ), .A1(n1046), .B0(\U4/U6/temp[3] ), .B1(
        n983), .Y(n1459) );
  AOI22X1 U1072 ( .A0(\U4/U6/temp[7] ), .A1(n1047), .B0(\U4/U6/temp[4] ), .B1(
        n986), .Y(n1460) );
  AOI2BB2X1 U1087 ( .B0(n2141), .B1(n1471), .A0N(n1471), .A1N(n2141), .Y(n1470) );
  MXI2X1 U1088 ( .A(n1463), .B(n968), .S0(n1472), .Y(\U4/Xt[5] ) );
  AOI2BB2X1 U1089 ( .B0(n1473), .B1(n1474), .A0N(n1473), .A1N(n1474), .Y(n1472) );
  MXI2X1 U1090 ( .A(n1463), .B(n968), .S0(n1475), .Y(\U4/Xt[4] ) );
  AOI2BB2X1 U1091 ( .B0(n1476), .B1(n1477), .A0N(n1477), .A1N(n1476), .Y(n1475) );
  AOI22X1 U1106 ( .A0(\U4/U5/temp[4] ), .A1(\U4/U5/temp[1] ), .B0(n1086), .B1(
        n1044), .Y(n1490) );
  AOI22X1 U1113 ( .A0(\U4/U5/temp[2] ), .A1(\U4/temp5t[2] ), .B0(n1066), .B1(
        n1087), .Y(n1495) );
  AOI2BB2X1 U1118 ( .B0(\U4/U5/temp[0] ), .B1(n1043), .A0N(n1043), .A1N(
        \U4/U5/temp[0] ), .Y(n1501) );
  AOI22X1 U1120 ( .A0(\U4/U5/temp[5] ), .A1(n1087), .B0(\U4/U5/temp[2] ), .B1(
        n1045), .Y(n1503) );
  AOI22X1 U1122 ( .A0(\U4/U5/temp[11] ), .A1(n971), .B0(\U4/U5/temp[6] ), .B1(
        n1019), .Y(n1504) );
  AOI2BB2X1 U1129 ( .B0(\U4/temp5t[1] ), .B1(n1086), .A0N(n1086), .A1N(
        \U4/temp5t[1] ), .Y(n1508) );
  AOI22X1 U1133 ( .A0(\U4/U5/temp[6] ), .A1(n1043), .B0(\U4/U5/temp[3] ), .B1(
        n971), .Y(n1511) );
  AOI22X1 U1135 ( .A0(\U4/U5/temp[7] ), .A1(n1044), .B0(\U4/U5/temp[4] ), .B1(
        n974), .Y(n1512) );
  OAI21XL U1174 ( .A0(n2567), .A1(\U5/temp2[0] ), .B0(\U5/temp1[0] ), .Y(n1520) );
  AOI2BB2X1 U1325 ( .B0(n1657), .B1(n1658), .A0N(n1658), .A1N(n1657), .Y(n1656) );
  AOI22X1 U1347 ( .A0(n1683), .A1(n1684), .B0(n735), .B1(n763), .Y(n1682) );
  AOI22X1 U1350 ( .A0(n752), .A1(n748), .B0(n1687), .B1(n1688), .Y(n1685) );
  AOI22X1 U1484 ( .A0(n1672), .A1(n1817), .B0(n751), .B1(n725), .Y(
        \U2/temp_x[0] ) );
  AOI2BB2X1 U1569 ( .B0(n1877), .B1(n651), .A0N(n651), .A1N(n1877), .Y(n1876)
         );
  AOI2BB2X1 U1571 ( .B0(n1880), .B1(n1881), .A0N(n1880), .A1N(n1881), .Y(n1879) );
  AOI2BB2X1 U1656 ( .B0(n1983), .B1(n1984), .A0N(n1984), .A1N(n1983), .Y(n1982) );
  OAI2BB1X1 U1727 ( .A0N(n639), .A1N(n2031), .B0(n638), .Y(\U1/temp_xxx[0] )
         );
  DFFHQX4 \U4/U12/temp_reg[3]  ( .D(n819), .CK(clk), .Q(\U4/U6/temp[0] ) );
  DFFHQX4 \U5/U12/temp_reg[3]  ( .D(\U5/temp7[3] ), .CK(clk), .Q(
        \U5/U6/temp[0] ) );
  DFFHQX4 \U5/U11/temp_reg[3]  ( .D(n796), .CK(clk), .Q(\U5/U5/temp[0] ) );
  DFFHQX4 \U4/U11/temp_reg[3]  ( .D(\U4/temp5[3] ), .CK(clk), .Q(
        \U4/U5/temp[0] ) );
  DFFHQX4 \U7/temp_reg[1]  ( .D(temp1[1]), .CK(clk), .Q(temp1t[1]) );
  DFFHQX4 \U8/temp_reg[1]  ( .D(temp2[1]), .CK(clk), .Q(temp2t[1]) );
  DFFHQXL \U5/U13/temp_reg[11]  ( .D(\U5/Xt[11] ), .CK(clk), .Q(result5[11])
         );
  DFFHQXL \U1/U21/temp_reg[10]  ( .D(\U1/temp_yyy[10] ), .CK(clk), .Q(
        \U1/result6[2] ) );
  DFFHQXL \U2/U20/temp_reg[11]  ( .D(\U2/temp_x[11] ), .CK(clk), .Q(
        \U2/result1[11] ) );
  DFFHQXL \U2/U21/temp_reg[11]  ( .D(\U2/temp_y[11] ), .CK(clk), .Q(
        \U2/result2[11] ) );
  DFFHQXL \U1/U20/temp_reg[10]  ( .D(\U1/temp_xxx[10] ), .CK(clk), .Q(
        \U1/result5[2] ) );
  DFFHQX2 \U5/U12/temp_reg[5]  ( .D(\U5/temp7[5] ), .CK(clk), .Q(
        \U5/U6/temp[2] ) );
  DFFHQX2 \U4/U11/temp_reg[5]  ( .D(\U4/temp5[5] ), .CK(clk), .Q(
        \U4/U5/temp[2] ) );
  DFFHQX2 \U4/U11/temp_reg[0]  ( .D(\U4/temp5[0] ), .CK(clk), .Q(
        \U4/temp5t[0] ) );
  AOI22X1 U1574 ( .A0(n2482), .A1(n2549), .B0(n654), .B1(n1853), .Y(n1883) );
  DFFHQX1 \U10/temp_reg[4]  ( .D(temp4[4]), .CK(clk), .Q(temp4t[4]) );
  DFFHQX2 \U3/U21/temp_reg[11]  ( .D(\U3/temp10[11] ), .CK(clk), .Q(
        \U3/temp11[1] ) );
  DFFHQX2 \U9/temp_reg[2]  ( .D(temp3[2]), .CK(clk), .Q(temp3t[2]) );
  DFFHQXL \U4/U14/temp_reg[9]  ( .D(\U4/Yt[9] ), .CK(clk), .Q(result4[9]) );
  DFFHQX1 \U12/temp_reg[9]  ( .D(temp6[9]), .CK(clk), .Q(\U4/temp1[9] ) );
  DFFHQX1 \U11/temp_reg[9]  ( .D(temp5[9]), .CK(clk), .Q(\U5/temp1[9] ) );
  DFFHQX1 \U12/temp_reg[8]  ( .D(temp6[8]), .CK(clk), .Q(\U4/temp1[7] ) );
  DFFHQXL \U1/U21/temp_reg[9]  ( .D(\U1/temp_yyy[9] ), .CK(clk), .Q(
        \U1/result6[1] ) );
  DFFHQXL \U1/U20/temp_reg[9]  ( .D(\U1/temp_xxx[9] ), .CK(clk), .Q(
        \U1/result5[1] ) );
  DFFHQX1 \U7/temp_reg[2]  ( .D(temp1[2]), .CK(clk), .Q(temp1t[2]) );
  DFFHQX1 \U7/temp_reg[4]  ( .D(temp1[4]), .CK(clk), .Q(temp1t[4]) );
  DFFHQX1 \U5/U12/temp_reg[0]  ( .D(\U5/temp7[0] ), .CK(clk), .Q(
        \U5/temp7t[0] ) );
  DFFHQX2 \U14/temp_reg[1]  ( .D(temp8[1]), .CK(clk), .Q(\U5/temp2[0] ) );
  DFFHQX2 \U10/temp_reg[2]  ( .D(temp4[2]), .CK(clk), .Q(temp4t[2]) );
  DFFHQX2 \U8/temp_reg[2]  ( .D(temp2[2]), .CK(clk), .Q(temp2t[2]) );
  DFFHQX2 \U7/temp_reg[3]  ( .D(temp1[3]), .CK(clk), .Q(temp1t[3]) );
  DFFHQX2 \U4/U12/temp_reg[5]  ( .D(n817), .CK(clk), .Q(\U4/U6/temp[2] ) );
  DFFHQX2 \U5/U11/temp_reg[5]  ( .D(n794), .CK(clk), .Q(\U5/U5/temp[2] ) );
  DFFHQX1 \U5/U12/temp_reg[1]  ( .D(\U5/temp7[1] ), .CK(clk), .Q(
        \U5/temp7t[1] ) );
  INVX1 U513 ( .A(n1447), .Y(n1067) );
  INVX1 U535 ( .A(\U4/U6/temp[2] ), .Y(n1089) );
  INVX1 U537 ( .A(\U5/U5/temp[2] ), .Y(n1091) );
  INVX1 U523 ( .A(n1390), .Y(n1077) );
  INVX1 U533 ( .A(\U4/U5/temp[2] ), .Y(n1087) );
  INVX1 U225 ( .A(n2053), .Y(n784) );
  INVX1 U227 ( .A(\intadd_39/A[1] ), .Y(n786) );
  INVX1 U148 ( .A(\intadd_35/B[2] ), .Y(n707) );
  INVX1 U152 ( .A(\intadd_35/B[1] ), .Y(n711) );
  INVX1 U156 ( .A(\intadd_35/CI ), .Y(n715) );
  INVX1 U162 ( .A(\intadd_45/SUM[1] ), .Y(n721) );
  INVX1 U155 ( .A(n1228), .Y(n714) );
  INVX1 U164 ( .A(\intadd_45/SUM[0] ), .Y(n723) );
  INVX1 U518 ( .A(n1338), .Y(n1072) );
  INVX1 U539 ( .A(\U5/U6/temp[2] ), .Y(n1093) );
  INVX1 U31 ( .A(x2[7]), .Y(n590) );
  INVX1 U3 ( .A(x0[7]), .Y(n562) );
  INVX8 U168 ( .A(n1664), .Y(n727) );
  NAND3X1 U1533 ( .A(n1231), .B(\U2/result2[9] ), .C(n889), .Y(n1254) );
  INVX1 U550 ( .A(n1255), .Y(n1104) );
  INVX1 U554 ( .A(\U2/temp_yt[0] ), .Y(n1108) );
  INVX1 U552 ( .A(\U2/result2[0] ), .Y(n1106) );
  INVX1 U549 ( .A(n1261), .Y(n1103) );
  INVX1 U553 ( .A(\U2/temp_xt[0] ), .Y(n1107) );
  INVX1 U551 ( .A(\U2/result1[0] ), .Y(n1105) );
  INVX1 U315 ( .A(result5[8]), .Y(n873) );
  INVX1 U314 ( .A(result5[7]), .Y(n872) );
  INVX1 U313 ( .A(result5[6]), .Y(n871) );
  INVX1 U339 ( .A(result5[5]), .Y(n897) );
  INVX1 U338 ( .A(result5[4]), .Y(n896) );
  INVX1 U337 ( .A(result5[3]), .Y(n895) );
  INVX1 U358 ( .A(result5[2]), .Y(n916) );
  INVX1 U357 ( .A(result5[1]), .Y(n915) );
  INVX1 U320 ( .A(result6[8]), .Y(n878) );
  INVX1 U319 ( .A(result6[7]), .Y(n877) );
  INVX1 U318 ( .A(result6[6]), .Y(n876) );
  INVX1 U344 ( .A(result6[5]), .Y(n902) );
  INVX1 U343 ( .A(result6[4]), .Y(n901) );
  INVX1 U342 ( .A(result6[3]), .Y(n900) );
  INVX1 U361 ( .A(result6[2]), .Y(n919) );
  INVX1 U360 ( .A(result6[1]), .Y(n918) );
  INVX1 U349 ( .A(\U6/temp4t[3] ), .Y(n907) );
  INVX1 U348 ( .A(\U6/temp4t[2] ), .Y(n906) );
  INVX1 U363 ( .A(\U6/temp4t[1] ), .Y(n921) );
  MXI2X2 U1341 ( .A(n758), .B(n1673), .S0(n1674), .Y(n1658) );
  XNOR2X1 U1065 ( .A(n1455), .B(n1456), .Y(n1447) );
  XNOR2X1 U1049 ( .A(n1442), .B(n1443), .Y(n1435) );
  XNOR2X1 U1054 ( .A(n1448), .B(n1449), .Y(n1431) );
  XNOR2X1 U1056 ( .A(n1450), .B(n1451), .Y(n1425) );
  XOR2X1 U1675 ( .A(n1997), .B(n1998), .Y(n1996) );
  XNOR2X1 U1671 ( .A(n1992), .B(n1993), .Y(n1991) );
  XNOR2X1 U974 ( .A(n1393), .B(n1394), .Y(n1368) );
  OAI2BB2X2 U1590 ( .B0(n1892), .B1(n661), .A0N(n1892), .A1N(n661), .Y(n1877)
         );
  XNOR2X1 U1587 ( .A(n2164), .B(n1890), .Y(n1888) );
  XOR2X1 U1583 ( .A(n1886), .B(n1887), .Y(n1884) );
  OAI2BB2X2 U1582 ( .B0(n1884), .B1(n2550), .A0N(n1884), .A1N(n2550), .Y(n1874) );
  XNOR2X1 U1117 ( .A(n1500), .B(n1501), .Y(n1483) );
  INVX8 U407 ( .A(n1464), .Y(n965) );
  XNOR2X1 U1119 ( .A(n1502), .B(n1503), .Y(n1477) );
  XOR2X1 U1400 ( .A(n1673), .B(n1738), .Y(n1736) );
  OAI2BB2X2 U1399 ( .B0(n1736), .B1(n2531), .A0N(n1736), .A1N(n2531), .Y(n1703) );
  INVX8 U219 ( .A(n1243), .Y(n778) );
  CLKINVX3 U546 ( .A(\U5/temp2[3] ), .Y(n1100) );
  AOI222X4 U1172 ( .A0(\U5/temp1[1] ), .A1(\U5/temp2[1] ), .B0(\U5/temp1[1] ), 
        .B1(n1266), .C0(\U5/temp2[1] ), .C1(n1266), .Y(n1277) );
  CLKINVX3 U251 ( .A(\U5/temp1[0] ), .Y(n810) );
  ADDFX2 \intadd_39/U8  ( .A(n2053), .B(\intadd_39/B[2] ), .CI(\intadd_39/n8 ), 
        .CO(\intadd_39/n7 ), .S(\intadd_35/A[2] ) );
  ADDFX2 \intadd_39/U7  ( .A(n783), .B(\intadd_39/B[3] ), .CI(\intadd_39/n7 ), 
        .CO(\intadd_39/n6 ), .S(\intadd_33/A[0] ) );
  ADDFX2 \intadd_39/U6  ( .A(n2059), .B(\intadd_39/B[4] ), .CI(\intadd_39/n6 ), 
        .CO(\intadd_39/n5 ), .S(\intadd_33/A[1] ) );
  ADDFX2 \intadd_39/U5  ( .A(n781), .B(\intadd_39/B[5] ), .CI(\intadd_39/n5 ), 
        .CO(\intadd_39/n4 ), .S(\intadd_33/A[2] ) );
  ADDFX2 \intadd_39/U4  ( .A(n2055), .B(\intadd_39/B[6] ), .CI(\intadd_39/n4 ), 
        .CO(\intadd_39/n3 ), .S(\intadd_33/A[3] ) );
  ADDFX2 \intadd_39/U3  ( .A(n779), .B(\intadd_39/B[7] ), .CI(\intadd_39/n3 ), 
        .CO(\intadd_39/n2 ), .S(\intadd_33/A[4] ) );
  ADDFX2 \intadd_45/U8  ( .A(n2054), .B(\intadd_39/B[1] ), .CI(\intadd_45/n8 ), 
        .CO(\intadd_45/n7 ), .S(\intadd_45/SUM[2] ) );
  ADDFX2 \intadd_45/U7  ( .A(n782), .B(\intadd_39/B[2] ), .CI(\intadd_45/n7 ), 
        .CO(\intadd_45/n6 ), .S(\intadd_35/CI ) );
  ADDFX2 \intadd_45/U6  ( .A(n2058), .B(\intadd_39/B[3] ), .CI(\intadd_45/n6 ), 
        .CO(\intadd_45/n5 ), .S(\intadd_35/B[1] ) );
  ADDFX2 \intadd_45/U5  ( .A(n780), .B(\intadd_39/B[4] ), .CI(\intadd_45/n5 ), 
        .CO(\intadd_45/n4 ), .S(\intadd_35/B[2] ) );
  ADDFX2 \intadd_45/U4  ( .A(n2056), .B(\intadd_39/B[5] ), .CI(\intadd_45/n4 ), 
        .CO(\intadd_45/n3 ), .S(\intadd_35/B[3] ) );
  ADDFX2 \intadd_45/U3  ( .A(n777), .B(\intadd_39/B[6] ), .CI(\intadd_45/n3 ), 
        .CO(\intadd_45/n2 ), .S(\intadd_35/B[4] ) );
  CLKINVX3 U136 ( .A(\intadd_35/B[5] ), .Y(n695) );
  ADDFX2 \intadd_33/U11  ( .A(\intadd_33/A[0] ), .B(n714), .CI(n723), .CO(
        \intadd_33/n10 ), .S(\intadd_33/SUM[0] ) );
  ADDFX2 \intadd_33/U10  ( .A(\intadd_33/A[1] ), .B(n721), .CI(\intadd_33/n10 ), .CO(\intadd_33/n9 ), .S(\intadd_33/SUM[1] ) );
  ADDFX2 \intadd_33/U9  ( .A(\intadd_33/A[2] ), .B(n719), .CI(\intadd_33/n9 ), 
        .CO(\intadd_33/n8 ), .S(\intadd_33/SUM[2] ) );
  ADDFX2 \intadd_33/U8  ( .A(\intadd_33/A[3] ), .B(n715), .CI(\intadd_33/n8 ), 
        .CO(\intadd_33/n7 ), .S(\intadd_33/SUM[3] ) );
  ADDFX2 \intadd_33/U7  ( .A(\intadd_33/A[4] ), .B(n711), .CI(\intadd_33/n7 ), 
        .CO(\intadd_33/n6 ), .S(\intadd_33/SUM[4] ) );
  ADDFX2 \intadd_33/U6  ( .A(\intadd_33/A[5] ), .B(n707), .CI(\intadd_33/n6 ), 
        .CO(\intadd_33/n5 ), .S(\intadd_33/SUM[5] ) );
  ADDFX2 U908 ( .A(\intadd_33/A[6] ), .B(n703), .CI(\intadd_33/n5 ), .CO(
        \intadd_33/n4 ), .S(\intadd_33/SUM[6] ) );
  ADDFX2 U907 ( .A(n691), .B(n699), .CI(\intadd_33/n4 ), .CO(\intadd_33/n3 ), 
        .S(\intadd_33/SUM[7] ) );
  ADDFX2 \intadd_47/U5  ( .A(n1096), .B(\U5/temp1[5] ), .CI(\intadd_47/n5 ), 
        .CO(\intadd_47/n4 ), .S(\intadd_38/B[4] ) );
  ADDFX2 \intadd_47/U4  ( .A(n1060), .B(\U5/temp1[6] ), .CI(\intadd_47/n4 ), 
        .CO(\intadd_47/n3 ), .S(\intadd_38/B[5] ) );
  ADDFX2 \intadd_47/U3  ( .A(n1097), .B(\U5/temp1[7] ), .CI(\intadd_47/n3 ), 
        .CO(\intadd_47/n2 ), .S(\intadd_38/B[6] ) );
  ADDFX2 \intadd_47/U2  ( .A(\U5/temp1[9] ), .B(n1013), .CI(\intadd_47/n2 ), 
        .CO(\intadd_47/n1 ), .S(\intadd_38/B[7] ) );
  ADDFX2 \intadd_48/U7  ( .A(\U5/temp1[2] ), .B(\U5/temp2[3] ), .CI(
        \intadd_48/n7 ), .CO(\intadd_48/n6 ), .S(\intadd_42/A[2] ) );
  ADDFX2 \intadd_48/U5  ( .A(\U5/temp1[4] ), .B(\U5/temp2[5] ), .CI(
        \intadd_48/n5 ), .CO(\intadd_48/n4 ), .S(\intadd_38/A[1] ) );
  ADDFX2 \intadd_48/U4  ( .A(\U5/temp1[5] ), .B(\U5/temp2[6] ), .CI(
        \intadd_48/n4 ), .CO(\intadd_48/n3 ), .S(\intadd_38/A[2] ) );
  ADDFX2 \intadd_48/U3  ( .A(\U5/temp1[6] ), .B(\U5/temp2[7] ), .CI(
        \intadd_48/n3 ), .CO(\intadd_48/n2 ), .S(\intadd_38/A[3] ) );
  ADDFX2 \intadd_48/U2  ( .A(\U5/temp2[9] ), .B(\U5/temp1[7] ), .CI(
        \intadd_48/n2 ), .CO(\intadd_48/n1 ), .S(\intadd_38/A[4] ) );
  ADDFX2 \intadd_42/U4  ( .A(\intadd_42/B[6] ), .B(\intadd_38/A[3] ), .CI(
        \intadd_42/n4 ), .CO(\intadd_42/n3 ), .S(\U5/temp7[7] ) );
  ADDFX2 \intadd_42/U3  ( .A(\intadd_42/B[6] ), .B(\intadd_38/A[4] ), .CI(
        \intadd_42/n3 ), .CO(\intadd_42/n2 ), .S(\U5/temp7[8] ) );
  ADDFX2 \intadd_42/U2  ( .A(\intadd_42/B[6] ), .B(\intadd_38/A[5] ), .CI(
        \intadd_42/n2 ), .CO(\intadd_42/n1 ), .S(\U5/temp7[9] ) );
  ADDFX2 \intadd_35/U10  ( .A(\intadd_35/A[1] ), .B(\intadd_35/B[1] ), .CI(
        \intadd_35/n10 ), .CO(\intadd_35/n9 ), .S(\intadd_35/SUM[1] ) );
  ADDFX2 \intadd_35/U9  ( .A(\intadd_35/A[2] ), .B(\intadd_35/B[2] ), .CI(
        \intadd_35/n9 ), .CO(\intadd_35/n8 ), .S(\intadd_35/SUM[2] ) );
  ADDFX2 \intadd_35/U6  ( .A(\intadd_33/A[2] ), .B(\intadd_35/B[5] ), .CI(
        \intadd_35/n6 ), .CO(\intadd_35/n5 ), .S(\intadd_35/SUM[5] ) );
  ADDFX2 \intadd_35/U5  ( .A(\intadd_33/A[3] ), .B(n688), .CI(\intadd_35/n5 ), 
        .CO(\intadd_35/n4 ), .S(\intadd_35/SUM[6] ) );
  ADDFX2 \intadd_35/U4  ( .A(n690), .B(\intadd_33/A[4] ), .CI(\intadd_35/n4 ), 
        .CO(\intadd_35/n3 ), .S(\intadd_35/SUM[7] ) );
  AOI222X4 U894 ( .A0(\U5/U6/temp[6] ), .A1(n1022), .B0(\U5/U6/temp[6] ), .B1(
        n1332), .C0(n1022), .C1(n1332), .Y(n1330) );
  XNOR2X1 U911 ( .A(n1341), .B(n1342), .Y(n1316) );
  ADDFX2 \intadd_46/U7  ( .A(\U4/temp1[3] ), .B(\U4/temp2[2] ), .CI(
        \intadd_46/n7 ), .CO(\intadd_46/n6 ), .S(\intadd_37/B[2] ) );
  ADDFX2 \intadd_46/U5  ( .A(\U4/temp1[5] ), .B(\U4/temp2[4] ), .CI(
        \intadd_46/n5 ), .CO(\intadd_46/n4 ), .S(\intadd_37/B[4] ) );
  ADDFX2 \intadd_46/U4  ( .A(\U4/temp1[6] ), .B(\U4/temp2[5] ), .CI(
        \intadd_46/n4 ), .CO(\intadd_46/n3 ), .S(\intadd_37/B[5] ) );
  ADDFX2 \intadd_46/U3  ( .A(\U4/temp1[7] ), .B(\U4/temp2[6] ), .CI(
        \intadd_46/n3 ), .CO(\intadd_46/n2 ), .S(\intadd_37/B[6] ) );
  AOI222X4 U1013 ( .A0(\intadd_46/n1 ), .A1(n1114), .B0(\intadd_46/n1 ), .B1(
        n1119), .C0(n1114), .C1(n1119), .Y(\intadd_41/B[6] ) );
  INVX1 U505 ( .A(\U4/temp1[1] ), .Y(n1059) );
  ADDFX2 \intadd_50/U3  ( .A(n1016), .B(\U4/temp2[6] ), .CI(\intadd_50/n3 ), 
        .CO(\intadd_50/n2 ), .S(\intadd_41/A[5] ) );
  ADDFX2 \intadd_41/U4  ( .A(\intadd_41/B[6] ), .B(\intadd_41/A[6] ), .CI(
        \intadd_41/n4 ), .CO(\intadd_41/n3 ), .S(\intadd_41/SUM[6] ) );
  ADDFX2 \intadd_41/U3  ( .A(\intadd_41/B[6] ), .B(\intadd_41/A[7] ), .CI(
        \intadd_41/n3 ), .CO(\intadd_41/n2 ), .S(\intadd_41/SUM[7] ) );
  ADDFX2 \intadd_41/U2  ( .A(\intadd_41/B[6] ), .B(\intadd_41/A[8] ), .CI(
        \intadd_41/n2 ), .CO(\intadd_41/n1 ), .S(\intadd_41/SUM[8] ) );
  ADDFX2 \intadd_38/U4  ( .A(\intadd_38/A[6] ), .B(\intadd_38/B[6] ), .CI(
        \intadd_38/n4 ), .CO(\intadd_38/n3 ), .S(\intadd_38/SUM[6] ) );
  ADDFX2 \intadd_38/U3  ( .A(\intadd_38/A[6] ), .B(\intadd_38/B[7] ), .CI(
        \intadd_38/n3 ), .CO(\intadd_38/n2 ), .S(\intadd_38/SUM[7] ) );
  ADDFX2 \intadd_38/U2  ( .A(\intadd_38/A[6] ), .B(n2060), .CI(\intadd_38/n2 ), 
        .CO(\intadd_38/n1 ), .S(\intadd_38/SUM[8] ) );
  ADDFX2 \intadd_25/U13  ( .A(\U1/result5[1] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n13 ), .CO(\intadd_25/n12 ), .S(\intadd_25/SUM[8] ) );
  ADDFX2 \intadd_25/U12  ( .A(\U1/result5[2] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n12 ), .CO(\intadd_25/SUM[10] ), .S(\intadd_25/SUM[9] ) );
  ADDFX2 \intadd_25/U6  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[6] ), .CI(
        \intadd_25/n6 ), .CO(\intadd_25/n5 ), .S(\U1/Xtt[6] ) );
  ADDFX2 \intadd_25/U5  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[7] ), .CI(
        \intadd_25/n5 ), .CO(\intadd_25/n4 ), .S(\U1/Xtt[7] ) );
  ADDFX2 \intadd_25/U4  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[8] ), .CI(
        \intadd_25/n4 ), .CO(\intadd_25/n3 ), .S(\U1/Xtt[8] ) );
  ADDFX2 \intadd_25/U3  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[9] ), .CI(
        \intadd_25/n3 ), .CO(\intadd_25/n2 ), .S(\U1/Xtt[9] ) );
  ADDFX2 \intadd_25/U2  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[10] ), .CI(
        \intadd_25/n2 ), .CO(\U1/Xtt[11] ), .S(\U1/Xtt[10] ) );
  ADDFX2 \intadd_26/U13  ( .A(\U1/result6[1] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n13 ), .CO(\intadd_26/n12 ), .S(\intadd_26/SUM[8] ) );
  ADDFX2 \intadd_26/U6  ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[6] ), .CI(
        \intadd_26/n6 ), .CO(\intadd_26/n5 ), .S(\U1/Ytt[6] ) );
  ADDFX2 \intadd_26/U5  ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[7] ), .CI(
        \intadd_26/n5 ), .CO(\intadd_26/n4 ), .S(\U1/Ytt[7] ) );
  ADDFX2 \intadd_26/U4  ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[8] ), .CI(
        \intadd_26/n4 ), .CO(\intadd_26/n3 ), .S(\U1/Ytt[8] ) );
  ADDFX2 \intadd_37/U5  ( .A(n823), .B(\intadd_37/B[5] ), .CI(\intadd_37/n5 ), 
        .CO(\intadd_37/n4 ), .S(\U4/temp5[6] ) );
  ADDFX2 \intadd_37/U4  ( .A(\intadd_37/A[6] ), .B(\intadd_37/B[6] ), .CI(
        \intadd_37/n4 ), .CO(\intadd_37/n3 ), .S(\U4/temp5[7] ) );
  ADDFX2 \intadd_37/U3  ( .A(\intadd_37/A[6] ), .B(\intadd_37/B[7] ), .CI(
        \intadd_37/n3 ), .CO(\intadd_37/n2 ), .S(\U4/temp5[8] ) );
  ADDFX2 \intadd_37/U2  ( .A(\intadd_37/A[6] ), .B(\intadd_37/B[8] ), .CI(
        \intadd_37/n2 ), .CO(\intadd_37/n1 ), .S(\U4/temp5[9] ) );
  AOI222X4 U608 ( .A0(x2[6]), .A1(n623), .B0(x2[6]), .B1(n593), .C0(n623), 
        .C1(n593), .Y(n1160) );
  AOI222X4 U576 ( .A0(x0[6]), .A1(n633), .B0(x0[6]), .B1(n565), .C0(n633), 
        .C1(n565), .Y(n1128) );
  XOR2X1 U839 ( .A(n1112), .B(n1286), .Y(\U6/temp3[9] ) );
  INVX1 U377 ( .A(\U4/temp2[7] ), .Y(n935) );
  INVX1 U466 ( .A(\U4/temp2[6] ), .Y(n1023) );
  INVX1 U467 ( .A(\U4/temp2[5] ), .Y(n1024) );
  INVX1 U458 ( .A(\U4/temp2[4] ), .Y(n1015) );
  INVX1 U457 ( .A(\U4/temp2[3] ), .Y(n1014) );
  INVX1 U502 ( .A(\U4/temp2[1] ), .Y(n1057) );
  INVX1 U354 ( .A(\U6/temp6[4] ), .Y(n912) );
  INVX1 U353 ( .A(\U6/temp6[3] ), .Y(n911) );
  INVX1 U352 ( .A(\U6/temp6[2] ), .Y(n910) );
  INVX1 U371 ( .A(\U6/temp6[1] ), .Y(n929) );
  XNOR2X1 U1014 ( .A(\intadd_41/A[2] ), .B(n1283), .Y(\U4/temp5[0] ) );
  XNOR2X1 U851 ( .A(\intadd_38/B[2] ), .B(n1262), .Y(\U5/temp7[0] ) );
  INVX8 U531 ( .A(temp4t[3]), .Y(n1085) );
  INVX8 U534 ( .A(\U4/U6/temp[1] ), .Y(n1088) );
  INVX1 U425 ( .A(\U4/U6/temp[6] ), .Y(n983) );
  XNOR2X1 U1042 ( .A(n1437), .B(n1438), .Y(n1428) );
  INVX8 U536 ( .A(\U5/U5/temp[1] ), .Y(n1090) );
  XNOR2X1 U983 ( .A(n1398), .B(n1399), .Y(n1390) );
  XOR2X2 U987 ( .A(n1401), .B(n1402), .Y(n1364) );
  XNOR2X1 U967 ( .A(n1385), .B(n1386), .Y(n1378) );
  XOR2X2 U1132 ( .A(n1510), .B(n1511), .Y(n1473) );
  XNOR2X1 U1128 ( .A(n1507), .B(n1508), .Y(n1499) );
  XNOR2X1 U1112 ( .A(n1494), .B(n1495), .Y(n1487) );
  OAI22X1 U803 ( .A0(n1097), .A1(n1115), .B0(\U5/temp1[6] ), .B1(\U5/temp2[6] ), .Y(n1246) );
  OAI22X1 U813 ( .A0(n1094), .A1(n1060), .B0(\U5/temp2[5] ), .B1(\U5/temp1[5] ), .Y(n1273) );
  OAI2BB2X1 U806 ( .B0(\U5/temp1[4] ), .B1(\U5/temp2[4] ), .A0N(\U5/temp2[4] ), 
        .A1N(\U5/temp1[4] ), .Y(n1248) );
  OAI22X1 U815 ( .A0(n1111), .A1(n1100), .B0(\U5/temp2[3] ), .B1(\U5/temp1[3] ), .Y(n1276) );
  INVX1 U224 ( .A(n2054), .Y(n783) );
  OAI2BB2X1 U809 ( .B0(\U5/temp1[2] ), .B1(\U5/temp2[2] ), .A0N(\U5/temp2[2] ), 
        .A1N(\U5/temp1[2] ), .Y(n1249) );
  INVX1 U223 ( .A(n2059), .Y(n782) );
  INVX1 U144 ( .A(\intadd_35/B[3] ), .Y(n703) );
  ADDFX2 \intadd_47/U7  ( .A(n1125), .B(\U5/temp1[3] ), .CI(\intadd_47/n7 ), 
        .CO(\intadd_47/n6 ), .S(\intadd_38/B[2] ) );
  INVX1 U243 ( .A(n2060), .Y(n802) );
  AOI21X1 U852 ( .A0(n800), .A1(n852), .B0(\intadd_48/CI ), .Y(n1262) );
  NOR2BX1 U794 ( .AN(n1262), .B(\intadd_38/B[2] ), .Y(\intadd_42/A[0] ) );
  INVX8 U538 ( .A(\U5/U6/temp[1] ), .Y(n1092) );
  XNOR2X1 U909 ( .A(n1339), .B(n1340), .Y(n1322) );
  XNOR2X1 U920 ( .A(n1346), .B(n1347), .Y(n1338) );
  XNOR2X1 U897 ( .A(n1333), .B(n1334), .Y(n1326) );
  XNOR2X1 U890 ( .A(n1328), .B(n1329), .Y(n1319) );
  INVX1 U331 ( .A(\U2/result2[11] ), .Y(n889) );
  AOI2BB2X1 U761 ( .B0(n1235), .B1(\U2/result2[5] ), .A0N(\U2/result2[5] ), 
        .A1N(n1235), .Y(n2065) );
  AOI21X1 U780 ( .A0(n937), .A1(n1253), .B0(n1235), .Y(\intadd_44/B[1] ) );
  AOI2BB2X1 U764 ( .B0(n1238), .B1(\U2/result2[3] ), .A0N(\U2/result2[3] ), 
        .A1N(n1238), .Y(n2068) );
  INVX1 U68 ( .A(x6[8]), .Y(n627) );
  INVX1 U16 ( .A(x1[8]), .Y(n575) );
  OAI22X1 U695 ( .A0(n627), .A1(n575), .B0(x1[8]), .B1(x6[8]), .Y(n1143) );
  INVX1 U376 ( .A(\U4/temp1[6] ), .Y(n934) );
  INVX1 U459 ( .A(\U4/temp1[5] ), .Y(n1016) );
  INVX1 U461 ( .A(\U4/temp1[4] ), .Y(n1018) );
  INVX1 U460 ( .A(\U4/temp1[3] ), .Y(n1017) );
  INVX1 U58 ( .A(x4[8]), .Y(n617) );
  INVX1 U44 ( .A(x3[8]), .Y(n603) );
  INVX1 U17 ( .A(x1[7]), .Y(n576) );
  INVX1 U69 ( .A(x6[6]), .Y(n628) );
  INVX1 U22 ( .A(x1[4]), .Y(n581) );
  INVX1 U45 ( .A(x3[7]), .Y(n604) );
  INVX1 U59 ( .A(x4[6]), .Y(n618) );
  INVX1 U50 ( .A(x3[4]), .Y(n609) );
  OAI22X1 U639 ( .A0(n617), .A1(n603), .B0(x3[8]), .B1(x4[8]), .Y(n1175) );
  NAND3X1 U1544 ( .A(n1232), .B(\U2/result1[9] ), .C(n888), .Y(n1260) );
  AOI21X1 U786 ( .A0(n913), .A1(n1257), .B0(n1232), .Y(\intadd_43/B[5] ) );
  AOI2BB2X1 U760 ( .B0(n1234), .B1(\U2/result1[7] ), .A0N(\U2/result1[7] ), 
        .A1N(n1234), .Y(n2064) );
  AOI21X1 U787 ( .A0(n930), .A1(n1258), .B0(n1234), .Y(\intadd_43/B[3] ) );
  AOI2BB2X1 U762 ( .B0(n1236), .B1(\U2/result1[5] ), .A0N(\U2/result1[5] ), 
        .A1N(n1236), .Y(n2066) );
  AOI21X1 U788 ( .A0(n936), .A1(n1259), .B0(n1236), .Y(\intadd_43/B[1] ) );
  AOI2BB2X1 U763 ( .B0(n1237), .B1(\U2/result1[3] ), .A0N(\U2/result1[3] ), 
        .A1N(n1237), .Y(n2067) );
  XNOR2X1 U1543 ( .A(\intadd_43/n1 ), .B(n1260), .Y(\U2/Xtt[9] ) );
  AOI2BB2X1 U642 ( .B0(x4[7]), .B1(x3[7]), .A0N(x3[7]), .A1N(x4[7]), .Y(n1177)
         );
  AOI2BB2X1 U623 ( .B0(n1177), .B1(n1176), .A0N(n1176), .A1N(n1177), .Y(
        temp5[7]) );
  AOI2BB2X1 U698 ( .B0(x6[7]), .B1(x1[7]), .A0N(x1[7]), .A1N(x6[7]), .Y(n1145)
         );
  AOI2BB2X1 U591 ( .B0(n1145), .B1(n1144), .A0N(n1144), .A1N(n1145), .Y(
        temp7[7]) );
  INVX1 U269 ( .A(\intadd_41/A[5] ), .Y(n827) );
  AOI21X1 U1015 ( .A0(n850), .A1(n1110), .B0(\intadd_46/CI ), .Y(n1283) );
  NOR2BX1 U822 ( .AN(n1283), .B(\intadd_41/A[2] ), .Y(\intadd_37/B[0] ) );
  INVX1 U64 ( .A(x5[6]), .Y(n623) );
  INVX1 U36 ( .A(x2[4]), .Y(n595) );
  INVX1 U66 ( .A(x5[3]), .Y(n625) );
  INVX1 U74 ( .A(x7[6]), .Y(n633) );
  INVX1 U8 ( .A(x0[4]), .Y(n567) );
  INVX1 U76 ( .A(x7[3]), .Y(n635) );
  INVX1 U63 ( .A(x5[8]), .Y(n622) );
  OAI22X1 U667 ( .A0(n622), .A1(n589), .B0(x2[8]), .B1(x5[8]), .Y(n1159) );
  AOI2BB2X1 U605 ( .B0(n1159), .B1(n1158), .A0N(n1158), .A1N(n1159), .Y(
        temp6[8]) );
  INVX1 U73 ( .A(x7[8]), .Y(n632) );
  OAI22X1 U723 ( .A0(n632), .A1(n561), .B0(x0[8]), .B1(x7[8]), .Y(n1127) );
  AOI2BB2X1 U573 ( .B0(n1127), .B1(n1126), .A0N(n1126), .A1N(n1127), .Y(
        temp8[8]) );
  MXI2X1 U697 ( .A(n1210), .B(n578), .S0(n1145), .Y(temp2[7]) );
  MXI2X1 U641 ( .A(n1192), .B(n606), .S0(n1177), .Y(temp4[7]) );
  AOI2BB2X1 U701 ( .B0(x1[6]), .B1(x6[6]), .A0N(x6[6]), .A1N(x1[6]), .Y(n1147)
         );
  AOI2BB2X1 U593 ( .B0(n1146), .B1(n1147), .A0N(n1147), .A1N(n1146), .Y(
        temp7[6]) );
  AOI2BB2X1 U645 ( .B0(x3[6]), .B1(x4[6]), .A0N(x4[6]), .A1N(x3[6]), .Y(n1179)
         );
  AOI2BB2X1 U625 ( .B0(n1178), .B1(n1179), .A0N(n1179), .A1N(n1178), .Y(
        temp5[6]) );
  MXI2X1 U700 ( .A(n1211), .B(n580), .S0(n1147), .Y(temp2[6]) );
  MXI2X1 U644 ( .A(n1193), .B(n608), .S0(n1179), .Y(temp4[6]) );
  AOI2BB2X1 U670 ( .B0(x5[7]), .B1(x2[7]), .A0N(x2[7]), .A1N(x5[7]), .Y(n1161)
         );
  AOI2BB2X1 U607 ( .B0(n1161), .B1(n1160), .A0N(n1160), .A1N(n1161), .Y(
        temp6[7]) );
  AOI2BB2X1 U726 ( .B0(x7[7]), .B1(x0[7]), .A0N(x0[7]), .A1N(x7[7]), .Y(n1129)
         );
  AOI2BB2X1 U575 ( .B0(n1129), .B1(n1128), .A0N(n1128), .A1N(n1129), .Y(
        temp8[7]) );
  MXI2X1 U669 ( .A(n1201), .B(n592), .S0(n1161), .Y(temp3[7]) );
  MXI2X1 U725 ( .A(n1219), .B(n564), .S0(n1129), .Y(temp1[7]) );
  OAI2BB2X1 U704 ( .B0(x1[5]), .B1(x6[5]), .A0N(x6[5]), .A1N(x1[5]), .Y(n1149)
         );
  MXI2X1 U703 ( .A(n582), .B(n1212), .S0(n1149), .Y(temp2[5]) );
  OAI2BB2X1 U648 ( .B0(x3[5]), .B1(x4[5]), .A0N(x4[5]), .A1N(x3[5]), .Y(n1181)
         );
  AOI2BB2X1 U627 ( .B0(n1180), .B1(n1181), .A0N(n1181), .A1N(n1180), .Y(
        temp5[5]) );
  AOI2BB2X1 U595 ( .B0(n1148), .B1(n1149), .A0N(n1149), .A1N(n1148), .Y(
        temp7[5]) );
  MXI2X1 U647 ( .A(n610), .B(n1194), .S0(n1181), .Y(temp4[5]) );
  INVX1 U159 ( .A(\intadd_35/B[0] ), .Y(n718) );
  AOI21X1 U752 ( .A0(\intadd_35/A[2] ), .A1(n765), .B0(n1228), .Y(n2049) );
  AOI2BB2X1 U729 ( .B0(x0[6]), .B1(x7[6]), .A0N(x7[6]), .A1N(x0[6]), .Y(n1131)
         );
  AOI2BB2X1 U577 ( .B0(n1130), .B1(n1131), .A0N(n1131), .A1N(n1130), .Y(
        temp8[6]) );
  AOI2BB2X1 U673 ( .B0(x2[6]), .B1(x5[6]), .A0N(x5[6]), .A1N(x2[6]), .Y(n1163)
         );
  AOI2BB2X1 U609 ( .B0(n1162), .B1(n1163), .A0N(n1163), .A1N(n1162), .Y(
        temp6[6]) );
  AOI2BB2X1 U707 ( .B0(x1[4]), .B1(x6[4]), .A0N(x6[4]), .A1N(x1[4]), .Y(n1151)
         );
  AOI2BB2X1 U597 ( .B0(n1150), .B1(n1151), .A0N(n1151), .A1N(n1150), .Y(
        temp7[4]) );
  AOI2BB2X1 U651 ( .B0(x3[4]), .B1(x4[4]), .A0N(x4[4]), .A1N(x3[4]), .Y(n1183)
         );
  AOI2BB2X1 U629 ( .B0(n1182), .B1(n1183), .A0N(n1183), .A1N(n1182), .Y(
        temp5[4]) );
  MXI2X1 U650 ( .A(n1195), .B(n611), .S0(n1183), .Y(temp4[4]) );
  INVX1 U236 ( .A(\intadd_38/SUM[3] ), .Y(n795) );
  MXI2X1 U672 ( .A(n1202), .B(n594), .S0(n1163), .Y(temp3[6]) );
  MXI2X1 U728 ( .A(n1220), .B(n566), .S0(n1131), .Y(temp1[6]) );
  OAI2BB2X1 U710 ( .B0(x1[3]), .B1(x6[3]), .A0N(x6[3]), .A1N(x1[3]), .Y(n1153)
         );
  AOI2BB2X1 U599 ( .B0(n1152), .B1(n1153), .A0N(n1153), .A1N(n1152), .Y(
        temp7[3]) );
  OAI2BB2X1 U654 ( .B0(x3[3]), .B1(x4[3]), .A0N(x4[3]), .A1N(x3[3]), .Y(n1185)
         );
  AOI2BB2X1 U631 ( .B0(n1184), .B1(n1185), .A0N(n1185), .A1N(n1184), .Y(
        temp5[3]) );
  AOI2BB2X1 U1064 ( .B0(n2543), .B1(n1447), .A0N(n1447), .A1N(n2543), .Y(n1454) );
  INVX1 U237 ( .A(\intadd_38/SUM[2] ), .Y(n796) );
  INVX1 U262 ( .A(\intadd_41/SUM[1] ), .Y(n820) );
  INVX1 U238 ( .A(\intadd_38/SUM[1] ), .Y(n797) );
  INVX1 U263 ( .A(\intadd_41/SUM[0] ), .Y(n821) );
  INVX1 U239 ( .A(\intadd_38/SUM[0] ), .Y(n798) );
  OAI21XL U1001 ( .A0(\intadd_37/B[2] ), .A1(n1406), .B0(n1407), .Y(
        \U4/temp7[0] ) );
  INVX1 U281 ( .A(\intadd_40/SUM[8] ), .Y(n839) );
  MXI2X1 U706 ( .A(n1213), .B(n583), .S0(n1151), .Y(temp2[4]) );
  INVX1 U298 ( .A(result2[11]), .Y(n856) );
  INVX1 U310 ( .A(result4[11]), .Y(n868) );
  INVX1 U297 ( .A(\intadd_30/n1 ), .Y(n855) );
  INVX1 U296 ( .A(result1[11]), .Y(n854) );
  INVX1 U309 ( .A(result3[11]), .Y(n867) );
  INVX1 U295 ( .A(\intadd_29/n1 ), .Y(n853) );
  INVX1 U305 ( .A(result7[11]), .Y(n863) );
  INVX1 U301 ( .A(result5[9]), .Y(n859) );
  INVX1 U299 ( .A(\intadd_31/SUM[9] ), .Y(n857) );
  INVX1 U306 ( .A(result8[11]), .Y(n864) );
  INVX1 U304 ( .A(result6[9]), .Y(n862) );
  INVX1 U302 ( .A(\intadd_32/SUM[9] ), .Y(n860) );
  INVX1 U282 ( .A(\intadd_40/SUM[7] ), .Y(n840) );
  OAI2BB2X1 U676 ( .B0(x2[5]), .B1(x5[5]), .A0N(x5[5]), .A1N(x2[5]), .Y(n1165)
         );
  AOI2BB2X1 U611 ( .B0(n1164), .B1(n1165), .A0N(n1165), .A1N(n1164), .Y(
        temp6[5]) );
  OAI2BB2X1 U732 ( .B0(x0[5]), .B1(x7[5]), .A0N(x7[5]), .A1N(x0[5]), .Y(n1133)
         );
  AOI2BB2X1 U579 ( .B0(n1132), .B1(n1133), .A0N(n1133), .A1N(n1132), .Y(
        temp8[5]) );
  INVX1 U300 ( .A(\intadd_31/SUM[8] ), .Y(n858) );
  INVX1 U303 ( .A(\intadd_32/SUM[8] ), .Y(n861) );
  INVX1 U333 ( .A(\U6/temp6[5] ), .Y(n891) );
  INVX1 U327 ( .A(\U6/temp5[10] ), .Y(n885) );
  INVX1 U368 ( .A(\U6/temp6[0] ), .Y(n926) );
  INVX1 U321 ( .A(\intadd_36/SUM[9] ), .Y(n879) );
  MXI2X1 U653 ( .A(n613), .B(n1196), .S0(n1185), .Y(temp4[3]) );
  OAI21XL U861 ( .A0(\intadd_47/CI ), .A1(n1299), .B0(n799), .Y(n1298) );
  NAND2BX1 U860 ( .AN(\intadd_38/B[0] ), .B(n1298), .Y(\U5/temp5[0] ) );
  INVX1 U283 ( .A(\intadd_40/SUM[6] ), .Y(n841) );
  INVX1 U566 ( .A(\U6/temp6[10] ), .Y(n1120) );
  INVX1 U326 ( .A(\intadd_34/n1 ), .Y(n884) );
  MXI2X1 U675 ( .A(n596), .B(n1203), .S0(n1165), .Y(temp3[5]) );
  MXI2X1 U731 ( .A(n568), .B(n1221), .S0(n1133), .Y(temp1[5]) );
  INVX1 U322 ( .A(\intadd_36/SUM[8] ), .Y(n880) );
  INVX1 U307 ( .A(\intadd_31/SUM[7] ), .Y(n865) );
  INVX1 U308 ( .A(\intadd_32/SUM[7] ), .Y(n866) );
  INVX1 U284 ( .A(\intadd_40/SUM[5] ), .Y(n842) );
  INVX1 U323 ( .A(\intadd_36/SUM[7] ), .Y(n881) );
  INVX1 U311 ( .A(\intadd_31/SUM[6] ), .Y(n869) );
  INVX1 U316 ( .A(\intadd_32/SUM[6] ), .Y(n874) );
  INVX1 U285 ( .A(\intadd_40/SUM[4] ), .Y(n843) );
  AOI2BB2X1 U713 ( .B0(x1[2]), .B1(x6[2]), .A0N(x6[2]), .A1N(x1[2]), .Y(n1155)
         );
  AOI2BB2X1 U601 ( .B0(n1154), .B1(n1155), .A0N(n1155), .A1N(n1154), .Y(
        temp7[2]) );
  AOI2BB2X1 U657 ( .B0(x3[2]), .B1(x4[2]), .A0N(x4[2]), .A1N(x3[2]), .Y(n1187)
         );
  AOI2BB2X1 U633 ( .B0(n1186), .B1(n1187), .A0N(n1187), .A1N(n1186), .Y(
        temp5[2]) );
  AOI2BB2X1 U735 ( .B0(x0[4]), .B1(x7[4]), .A0N(x7[4]), .A1N(x0[4]), .Y(n1135)
         );
  MXI2X1 U734 ( .A(n1222), .B(n569), .S0(n1135), .Y(temp1[4]) );
  AOI2BB2X1 U679 ( .B0(x2[4]), .B1(x5[4]), .A0N(x5[4]), .A1N(x2[4]), .Y(n1167)
         );
  MXI2X1 U678 ( .A(n1204), .B(n597), .S0(n1167), .Y(temp3[4]) );
  INVX1 U324 ( .A(\intadd_36/SUM[6] ), .Y(n882) );
  INVX1 U317 ( .A(\intadd_32/SUM[5] ), .Y(n875) );
  INVX1 U312 ( .A(\intadd_31/SUM[5] ), .Y(n870) );
  INVX1 U286 ( .A(\intadd_40/SUM[3] ), .Y(n844) );
  MXI2X1 U709 ( .A(n585), .B(n1214), .S0(n1153), .Y(temp2[3]) );
  INVX1 U325 ( .A(\intadd_36/SUM[5] ), .Y(n883) );
  INVX1 U328 ( .A(\intadd_31/SUM[4] ), .Y(n886) );
  INVX1 U329 ( .A(\intadd_32/SUM[4] ), .Y(n887) );
  INVX1 U287 ( .A(\intadd_40/SUM[2] ), .Y(n845) );
  INVX1 U332 ( .A(\intadd_36/SUM[4] ), .Y(n890) );
  INVX1 U335 ( .A(\intadd_31/SUM[3] ), .Y(n893) );
  INVX1 U340 ( .A(\intadd_32/SUM[3] ), .Y(n898) );
  INVX1 U288 ( .A(\intadd_40/SUM[1] ), .Y(n846) );
  MXI2X1 U656 ( .A(n1197), .B(n614), .S0(n1187), .Y(temp4[2]) );
  MXI2X1 U712 ( .A(n1215), .B(n586), .S0(n1155), .Y(temp2[2]) );
  INVX1 U289 ( .A(\intadd_40/SUM[0] ), .Y(n847) );
  INVX1 U345 ( .A(\intadd_36/SUM[3] ), .Y(n903) );
  INVX1 U341 ( .A(\intadd_32/SUM[2] ), .Y(n899) );
  INVX1 U336 ( .A(\intadd_31/SUM[2] ), .Y(n894) );
  AOI2BB2X1 U613 ( .B0(n1166), .B1(n1167), .A0N(n1167), .A1N(n1166), .Y(
        temp6[4]) );
  AOI2BB2X1 U581 ( .B0(n1134), .B1(n1135), .A0N(n1135), .A1N(n1134), .Y(
        temp8[4]) );
  INVX1 U346 ( .A(\intadd_36/SUM[2] ), .Y(n904) );
  OAI2BB2X1 U738 ( .B0(x0[3]), .B1(x7[3]), .A0N(x7[3]), .A1N(x0[3]), .Y(n1137)
         );
  MXI2X1 U737 ( .A(n571), .B(n1223), .S0(n1137), .Y(temp1[3]) );
  OAI2BB2X1 U682 ( .B0(x2[3]), .B1(x5[3]), .A0N(x5[3]), .A1N(x2[3]), .Y(n1169)
         );
  MXI2X1 U681 ( .A(n599), .B(n1205), .S0(n1169), .Y(temp3[3]) );
  INVX1 U350 ( .A(\intadd_31/SUM[1] ), .Y(n908) );
  INVX1 U351 ( .A(\intadd_32/SUM[1] ), .Y(n909) );
  INVX1 U347 ( .A(\intadd_36/SUM[1] ), .Y(n905) );
  OAI2BB2X1 U688 ( .B0(x5[1]), .B1(x2[1]), .A0N(x2[1]), .A1N(x5[1]), .Y(n1173)
         );
  MXI2X1 U687 ( .A(n601), .B(n1207), .S0(n1173), .Y(temp3[1]) );
  AOI2BB2X1 U685 ( .B0(x2[2]), .B1(x5[2]), .A0N(x5[2]), .A1N(x2[2]), .Y(n1171)
         );
  MXI2X1 U684 ( .A(n1206), .B(n600), .S0(n1171), .Y(temp3[2]) );
  AOI2BB2X1 U741 ( .B0(x0[2]), .B1(x7[2]), .A0N(x7[2]), .A1N(x0[2]), .Y(n1139)
         );
  MXI2X1 U740 ( .A(n1224), .B(n572), .S0(n1139), .Y(temp1[2]) );
  OAI2BB2X1 U744 ( .B0(x7[1]), .B1(x0[1]), .A0N(x0[1]), .A1N(x7[1]), .Y(n1141)
         );
  MXI2X1 U743 ( .A(n573), .B(n1225), .S0(n1141), .Y(temp1[1]) );
  OAI2BB2X1 U716 ( .B0(x6[1]), .B1(x1[1]), .A0N(x1[1]), .A1N(x6[1]), .Y(n1157)
         );
  MXI2X1 U715 ( .A(n587), .B(n1216), .S0(n1157), .Y(temp2[1]) );
  OAI2BB2X1 U660 ( .B0(x4[1]), .B1(x3[1]), .A0N(x3[1]), .A1N(x4[1]), .Y(n1189)
         );
  MXI2X1 U659 ( .A(n615), .B(n1198), .S0(n1189), .Y(temp4[1]) );
  INVX1 U359 ( .A(\intadd_32/SUM[0] ), .Y(n917) );
  INVX1 U356 ( .A(\intadd_31/SUM[0] ), .Y(n914) );
  AOI2BB2X1 U583 ( .B0(n1136), .B1(n1137), .A0N(n1137), .A1N(n1136), .Y(
        temp8[3]) );
  AOI2BB2X1 U615 ( .B0(n1168), .B1(n1169), .A0N(n1169), .A1N(n1168), .Y(
        temp6[3]) );
  INVX1 U362 ( .A(\intadd_36/SUM[0] ), .Y(n920) );
  AOI2BB2X1 U585 ( .B0(n1138), .B1(n1139), .A0N(n1139), .A1N(n1138), .Y(
        temp8[2]) );
  AOI2BB2X1 U617 ( .B0(n1170), .B1(n1171), .A0N(n1171), .A1N(n1170), .Y(
        temp6[2]) );
  INVX8 U169 ( .A(n2560), .Y(n728) );
  NOR3X4 U1430 ( .A(n1721), .B(n1713), .C(n2434), .Y(n1763) );
  INVX1 U492 ( .A(\U4/U6/temp[4] ), .Y(n1047) );
  CLKINVX3 U280 ( .A(n1951), .Y(n838) );
  XNOR2X1 U972 ( .A(n1391), .B(n1392), .Y(n1374) );
  XNOR2X1 U960 ( .A(n1380), .B(n1381), .Y(n1371) );
  INVX8 U429 ( .A(n1357), .Y(n987) );
  INVX4 U278 ( .A(n1930), .Y(n836) );
  OAI2BB2X1 U1586 ( .B0(n1888), .B1(n1886), .A0N(n1888), .A1N(n1886), .Y(n1880) );
  NAND2X1 U1164 ( .A(\U5/temp2[9] ), .B(\U5/temp1[9] ), .Y(n1295) );
  OAI22X1 U811 ( .A0(n1056), .A1(n1013), .B0(\U5/temp2[7] ), .B1(\U5/temp1[7] ), .Y(n1270) );
  NOR2X1 U772 ( .A(n1240), .B(\intadd_39/A[0] ), .Y(\intadd_45/CI ) );
  NOR2X1 U864 ( .A(n2541), .B(n810), .Y(\intadd_47/CI ) );
  NOR2X1 U853 ( .A(n800), .B(n852), .Y(\intadd_48/CI ) );
  AOI2BB2X1 U819 ( .B0(n1098), .B1(\intadd_48/n1 ), .A0N(\intadd_48/n1 ), 
        .A1N(n1098), .Y(\intadd_38/A[5] ) );
  AOI22X1 U793 ( .A0(n1098), .A1(n804), .B0(\intadd_47/n1 ), .B1(n1244), .Y(
        n2060) );
  INVX1 U246 ( .A(\intadd_38/B[7] ), .Y(n805) );
  INVX1 U247 ( .A(\intadd_38/B[6] ), .Y(n806) );
  INVX1 U248 ( .A(\intadd_38/B[5] ), .Y(n807) );
  INVX1 U250 ( .A(\intadd_38/B[3] ), .Y(n809) );
  INVX1 U498 ( .A(\U5/U6/temp[4] ), .Y(n1053) );
  INVX4 U448 ( .A(n1312), .Y(n1006) );
  XOR2X2 U892 ( .A(n1330), .B(n1331), .Y(n1303) );
  INVX1 U334 ( .A(\U2/result2[8] ), .Y(n892) );
  INVX1 U379 ( .A(\U2/result2[4] ), .Y(n937) );
  CLKINVX3 U27 ( .A(n1215), .Y(n586) );
  CLKINVX3 U26 ( .A(n1214), .Y(n585) );
  CLKINVX3 U23 ( .A(n1212), .Y(n582) );
  CLKINVX3 U21 ( .A(n1211), .Y(n580) );
  NOR2X1 U843 ( .A(n1287), .B(n1288), .Y(n1289) );
  ADDFX2 \intadd_46/U2  ( .A(\U4/temp1[9] ), .B(\U4/temp2[7] ), .CI(
        \intadd_46/n2 ), .CO(\intadd_46/n1 ), .S(\intadd_37/B[7] ) );
  INVX1 U71 ( .A(x6[3]), .Y(n630) );
  INVX1 U25 ( .A(x1[2]), .Y(n584) );
  INVX1 U72 ( .A(x6[1]), .Y(n631) );
  INVX1 U61 ( .A(x4[3]), .Y(n620) );
  INVX1 U53 ( .A(x3[2]), .Y(n612) );
  INVX1 U62 ( .A(x4[1]), .Y(n621) );
  AOI2BB2X1 U756 ( .B0(n1232), .B1(\U2/result1[9] ), .A0N(\U2/result1[9] ), 
        .A1N(n1232), .Y(n2062) );
  AOI21X1 U1545 ( .A0(n1232), .A1(\U2/result1[9] ), .B0(n888), .Y(\U2/Xtt[10] ) );
  INVX1 U268 ( .A(\intadd_41/A[6] ), .Y(n826) );
  INVX1 U270 ( .A(\intadd_41/A[4] ), .Y(n828) );
  INVX1 U271 ( .A(\intadd_41/A[3] ), .Y(n829) );
  INVX1 U30 ( .A(x2[8]), .Y(n589) );
  INVX1 U39 ( .A(x2[2]), .Y(n598) );
  INVX1 U67 ( .A(x5[1]), .Y(n626) );
  INVX1 U2 ( .A(x0[8]), .Y(n561) );
  INVX1 U11 ( .A(x0[2]), .Y(n570) );
  INVX1 U77 ( .A(x7[1]), .Y(n636) );
  INVX1 U232 ( .A(\intadd_38/SUM[6] ), .Y(n791) );
  INVX1 U231 ( .A(\intadd_38/SUM[7] ), .Y(n790) );
  INVX1 U230 ( .A(\intadd_38/SUM[8] ), .Y(n789) );
  INVX1 U255 ( .A(\intadd_41/SUM[7] ), .Y(n814) );
  INVX1 U256 ( .A(\intadd_41/SUM[6] ), .Y(n815) );
  AOI2BB2X1 U1030 ( .B0(n1427), .B1(n1428), .A0N(n1428), .A1N(n1427), .Y(n1426) );
  INVX1 U143 ( .A(\intadd_33/SUM[2] ), .Y(n702) );
  AOI2BB2X1 U1095 ( .B0(n1482), .B1(n1483), .A0N(n1483), .A1N(n1482), .Y(n1481) );
  AOI2BB2X1 U880 ( .B0(n1321), .B1(n1322), .A0N(n1322), .A1N(n1321), .Y(n1320)
         );
  INVX1 U147 ( .A(\intadd_33/SUM[1] ), .Y(n706) );
  INVX1 U153 ( .A(\intadd_35/SUM[1] ), .Y(n712) );
  INVX1 U157 ( .A(\intadd_35/SUM[0] ), .Y(n716) );
  INVX1 U151 ( .A(\intadd_33/SUM[0] ), .Y(n710) );
  INVX1 U257 ( .A(\intadd_41/SUM[5] ), .Y(n816) );
  INVX1 U233 ( .A(\intadd_38/SUM[5] ), .Y(n792) );
  AOI2BB2X1 U982 ( .B0(n1389), .B1(n1390), .A0N(n1390), .A1N(n1389), .Y(n1397)
         );
  AOI2BB2X1 U1127 ( .B0(n1498), .B1(n1499), .A0N(n1499), .A1N(n1498), .Y(n1506) );
  INVX1 U260 ( .A(\intadd_41/SUM[3] ), .Y(n818) );
  INVX1 U261 ( .A(\intadd_41/SUM[2] ), .Y(n819) );
  AOI2BB2X1 U919 ( .B0(n1337), .B1(n1338), .A0N(n1338), .A1N(n1337), .Y(n1345)
         );
  INVX4 U199 ( .A(n1673), .Y(n758) );
  CLKINVX3 U491 ( .A(\U4/U6/temp[3] ), .Y(n1046) );
  XNOR2X2 U976 ( .A(n1384), .B(n1395), .Y(n1358) );
  INVX1 U495 ( .A(\U5/U5/temp[4] ), .Y(n1050) );
  INVX8 U101 ( .A(n1911), .Y(n660) );
  INVX8 U412 ( .A(n1473), .Y(n970) );
  XNOR2X1 U1105 ( .A(n1489), .B(n1490), .Y(n1480) );
  XOR2X1 U1393 ( .A(n1687), .B(n1730), .Y(n1729) );
  AOI2BB2X1 U814 ( .B0(n1280), .B1(n1276), .A0N(n1276), .A1N(n1280), .Y(n2054)
         );
  AOI2BB2X1 U776 ( .B0(n785), .B1(n1249), .A0N(n1249), .A1N(n785), .Y(n2053)
         );
  MXI2X1 U808 ( .A(n720), .B(n1277), .S0(n1249), .Y(\intadd_39/B[1] ) );
  INVX1 U206 ( .A(n1239), .Y(n765) );
  AOI22X1 U857 ( .A0(n803), .A1(n793), .B0(\intadd_38/A[6] ), .B1(
        \intadd_42/B[6] ), .Y(n1292) );
  INVX1 U249 ( .A(\intadd_38/B[4] ), .Y(n808) );
  CLKINVX3 U497 ( .A(\U5/U6/temp[3] ), .Y(n1052) );
  NAND3X1 U1542 ( .A(\U2/temp_yt[0] ), .B(\U2/result2[0] ), .C(\U2/result2[1] ), .Y(n1255) );
  AOI21X1 U1534 ( .A0(n1231), .A1(\U2/result2[9] ), .B0(n889), .Y(\U2/Ytt[10] ) );
  NOR2X1 U1011 ( .A(\U4/temp2[9] ), .B(\U4/temp1[7] ), .Y(n1287) );
  AOI22X1 U1008 ( .A0(n848), .A1(n825), .B0(\intadd_37/A[6] ), .B1(
        \intadd_41/B[6] ), .Y(n1405) );
  AOI22X1 U841 ( .A0(\U4/temp2[9] ), .A1(\U4/temp1[9] ), .B0(n1119), .B1(n1114), .Y(n1263) );
  INVX1 U558 ( .A(n1263), .Y(n1112) );
  ADDFX2 \intadd_50/U2  ( .A(n934), .B(\U4/temp2[7] ), .CI(\intadd_50/n2 ), 
        .CO(\intadd_50/n1 ), .S(\intadd_41/A[6] ) );
  AOI2BB2X1 U821 ( .B0(\intadd_46/n1 ), .B1(n1263), .A0N(n1263), .A1N(
        \intadd_46/n1 ), .Y(\intadd_37/B[8] ) );
  INVX1 U240 ( .A(\intadd_42/A[2] ), .Y(n799) );
  NAND3X1 U1553 ( .A(\U2/temp_xt[0] ), .B(\U2/result1[0] ), .C(\U2/result1[1] ), .Y(n1261) );
  INVX1 U266 ( .A(\intadd_41/A[7] ), .Y(n824) );
  INVX1 U34 ( .A(n1162), .Y(n593) );
  INVX1 U6 ( .A(n1130), .Y(n565) );
  INVX1 U254 ( .A(\intadd_41/SUM[8] ), .Y(n813) );
  MXI2X1 U945 ( .A(n1354), .B(n992), .S0(n1366), .Y(\U5/Xt[4] ) );
  INVX1 U139 ( .A(\intadd_33/SUM[3] ), .Y(n698) );
  INVX1 U145 ( .A(\intadd_35/SUM[3] ), .Y(n704) );
  AOI2BB2X1 U950 ( .B0(n1373), .B1(n1374), .A0N(n1374), .A1N(n1373), .Y(n1372)
         );
  INVX1 U149 ( .A(\intadd_35/SUM[2] ), .Y(n708) );
  OAI21XL U753 ( .A0(\intadd_45/SUM[2] ), .A1(n1229), .B0(n718), .Y(n2051) );
  MXI2X1 U1126 ( .A(n2141), .B(n1488), .S0(n1506), .Y(\U4/Xt[0] ) );
  MXI2X1 U1063 ( .A(n984), .B(n1436), .S0(n1454), .Y(\U4/Yt[0] ) );
  OAI21XL U1348 ( .A0(n1685), .A1(n747), .B0(n2529), .Y(\U2/temp_y[0] ) );
  NOR2X1 U832 ( .A(n923), .B(n925), .Y(\intadd_30/CI ) );
  NOR2X1 U833 ( .A(n922), .B(n924), .Y(\intadd_29/CI ) );
  NAND2X1 U758 ( .A(result7[0]), .B(n932), .Y(n1227) );
  INVX1 U369 ( .A(n1227), .Y(n927) );
  NAND2X1 U759 ( .A(result8[0]), .B(n933), .Y(n1226) );
  INVX1 U370 ( .A(n1226), .Y(n928) );
  INVX1 U403 ( .A(temp2t[8]), .Y(n961) );
  AOI2BB2X1 U1724 ( .B0(temp2t[8]), .B1(temp3t[8]), .A0N(temp3t[8]), .A1N(
        temp2t[8]), .Y(n1810) );
  CLKINVX3 U494 ( .A(\U5/U5/temp[3] ), .Y(n1049) );
  INVX8 U430 ( .A(n1367), .Y(n988) );
  OAI21XL U1620 ( .A0(n752), .A1(n1893), .B0(n1890), .Y(n1933) );
  CLKINVX3 U488 ( .A(\U4/U5/temp[3] ), .Y(n1043) );
  INVX1 U192 ( .A(n1817), .Y(n751) );
  CLKINVX3 U557 ( .A(\U5/temp1[3] ), .Y(n1111) );
  AOI22X4 U773 ( .A0(n1243), .A1(n1244), .B0(n1098), .B1(n778), .Y(n2057) );
  NAND2X1 U717 ( .A(x1[0]), .B(x6[0]), .Y(n1216) );
  NAND2X1 U661 ( .A(x3[0]), .B(x4[0]), .Y(n1198) );
  INVX1 U20 ( .A(n1146), .Y(n579) );
  INVX1 U48 ( .A(n1178), .Y(n607) );
  INVX1 U265 ( .A(\intadd_41/A[8] ), .Y(n823) );
  INVX1 U43 ( .A(x2[0]), .Y(n602) );
  INVX1 U15 ( .A(x0[0]), .Y(n574) );
  MXI2X1 U1027 ( .A(n1411), .B(n980), .S0(n1423), .Y(\U4/Yt[4] ) );
  NAND2X1 U689 ( .A(x2[0]), .B(x5[0]), .Y(n1207) );
  NAND2X1 U745 ( .A(x0[0]), .B(x7[0]), .Y(n1225) );
  INVX1 U138 ( .A(\intadd_33/SUM[4] ), .Y(n697) );
  AOI2BB2X1 U948 ( .B0(n1370), .B1(n1371), .A0N(n1371), .A1N(n1370), .Y(n1369)
         );
  INVX1 U141 ( .A(\intadd_35/SUM[4] ), .Y(n700) );
  AOI2BB2X1 U878 ( .B0(n1318), .B1(n1319), .A0N(n1319), .A1N(n1318), .Y(n1317)
         );
  MXI2X1 U1031 ( .A(n2138), .B(n1415), .S0(n1429), .Y(\U4/Yt[2] ) );
  MXI2X1 U1570 ( .A(n1867), .B(n659), .S0(n1879), .Y(\U1/temp_yyy[1] ) );
  MXI2X1 U981 ( .A(n996), .B(n1379), .S0(n1397), .Y(\U5/Xt[0] ) );
  INVX1 U90 ( .A(n1932), .Y(n649) );
  AOI2BB2X1 U1327 ( .B0(n2529), .B1(n1662), .A0N(n1662), .A1N(n2529), .Y(n1660) );
  MXI2X1 U918 ( .A(n1008), .B(n1327), .S0(n1345), .Y(\U5/Yt[0] ) );
  INVX1 U365 ( .A(result4[0]), .Y(n923) );
  INVX1 U367 ( .A(result2[0]), .Y(n925) );
  INVX1 U364 ( .A(result3[0]), .Y(n922) );
  INVX1 U366 ( .A(result1[0]), .Y(n924) );
  INVX1 U374 ( .A(result5[0]), .Y(n932) );
  INVX1 U375 ( .A(result6[0]), .Y(n933) );
  INVX1 U402 ( .A(temp1t[8]), .Y(n960) );
  AOI2BB2X1 U1720 ( .B0(temp4t[8]), .B1(temp1t[8]), .A0N(temp1t[8]), .A1N(
        temp4t[8]), .Y(n1812) );
  MXI2X1 U1344 ( .A(n759), .B(n2146), .S0(n1678), .Y(n1662) );
  INVX1 U548 ( .A(\U2/result2[2] ), .Y(n1102) );
  NAND2X1 U1540 ( .A(n1238), .B(\U2/result2[3] ), .Y(n1253) );
  AOI2BB2X1 U797 ( .B0(\intadd_50/n1 ), .B1(n1113), .A0N(n1113), .A1N(
        \intadd_50/n1 ), .Y(\intadd_41/A[7] ) );
  INVX1 U29 ( .A(x1[0]), .Y(n588) );
  NAND2X1 U719 ( .A(n588), .B(x6[0]), .Y(n1156) );
  INVX1 U57 ( .A(x3[0]), .Y(n616) );
  NAND2X1 U663 ( .A(n616), .B(x4[0]), .Y(n1188) );
  INVX1 U547 ( .A(\U2/result1[2] ), .Y(n1101) );
  MXI2X1 U1086 ( .A(n1463), .B(n968), .S0(n1470), .Y(\U4/Xt[6] ) );
  AOI222X4 U606 ( .A0(x5[7]), .A1(n590), .B0(x5[7]), .B1(n1160), .C0(n590), 
        .C1(n1160), .Y(n1158) );
  AOI222X4 U574 ( .A0(x7[7]), .A1(n562), .B0(x7[7]), .B1(n1128), .C0(n562), 
        .C1(n1128), .Y(n1126) );
  AOI2BB2X1 U1093 ( .B0(n1479), .B1(n1480), .A0N(n1480), .A1N(n1479), .Y(n1478) );
  MXI2X1 U949 ( .A(n2139), .B(n1358), .S0(n1372), .Y(\U5/Xt[2] ) );
  MXI2X1 U1094 ( .A(n966), .B(n1467), .S0(n1481), .Y(\U4/Xt[2] ) );
  MXI2X1 U879 ( .A(n1002), .B(n1306), .S0(n1320), .Y(\U5/Yt[2] ) );
  AOI2BB2X1 U1366 ( .B0(n1705), .B1(n1706), .A0N(n1705), .A1N(n1706), .Y(n1704) );
  INVX1 U504 ( .A(\U4/temp2[2] ), .Y(n1058) );
  CLKINVX3 U483 ( .A(temp3t[5]), .Y(n1038) );
  AOI22X1 U1715 ( .A0(temp2t[7]), .A1(n1039), .B0(temp3t[7]), .B1(n1037), .Y(
        n1799) );
  INVX1 U489 ( .A(\U4/U5/temp[4] ), .Y(n1044) );
  OAI2BB2X1 U1397 ( .B0(n1734), .B1(n763), .A0N(n1734), .A1N(n763), .Y(n1705)
         );
  INVX1 U190 ( .A(n1707), .Y(n749) );
  INVX1 U561 ( .A(\U5/temp1[6] ), .Y(n1115) );
  INVX1 U507 ( .A(\U4/temp1[2] ), .Y(n1061) );
  OAI21XL U1010 ( .A0(\U4/temp1[9] ), .A1(n1287), .B0(\intadd_50/n1 ), .Y(
        n1408) );
  AOI2BB2X1 U1652 ( .B0(n2345), .B1(n1977), .A0N(n1977), .A1N(n2345), .Y(n1976) );
  MXI2X1 U1029 ( .A(n1412), .B(n977), .S0(n1426), .Y(\U4/Yt[3] ) );
  AOI2BB2X1 U1364 ( .B0(n1702), .B1(n1703), .A0N(n1702), .A1N(n1703), .Y(n1701) );
  MXI2X1 U1655 ( .A(n646), .B(n2554), .S0(n1982), .Y(\U1/temp_xxx[1] ) );
  CLKINVX3 U477 ( .A(temp2t[4]), .Y(n1034) );
  AOI2BB2X1 U1738 ( .B0(temp2t[6]), .B1(temp3t[6]), .A0N(temp3t[6]), .A1N(
        temp2t[6]), .Y(n1808) );
  OAI21XL U1729 ( .A0(n752), .A1(n676), .B0(n1993), .Y(n2031) );
  AOI2BB2X2 U775 ( .B0(n1247), .B1(n1248), .A0N(n1248), .A1N(n1247), .Y(n2059)
         );
  INVX1 U134 ( .A(\intadd_33/SUM[5] ), .Y(n693) );
  INVX1 U137 ( .A(\intadd_35/SUM[5] ), .Y(n696) );
  AOI2BB2X1 U1321 ( .B0(n1650), .B1(n725), .A0N(n725), .A1N(n1650), .Y(n1649)
         );
  MXI2X1 U947 ( .A(n1355), .B(n989), .S0(n1369), .Y(\U5/Xt[3] ) );
  MXI2X1 U877 ( .A(n1303), .B(n1001), .S0(n1317), .Y(\U5/Yt[3] ) );
  INVX1 U92 ( .A(n1878), .Y(n651) );
  MXI2X1 U1568 ( .A(n2552), .B(n658), .S0(n1876), .Y(\U1/temp_yyy[2] ) );
  AOI2BB2X1 U1654 ( .B0(n1980), .B1(n1981), .A0N(n1981), .A1N(n1980), .Y(n1979) );
  AOI2BB2X1 U1368 ( .B0(n1709), .B1(n2555), .A0N(n1709), .A1N(n2555), .Y(n1708) );
  MXI2X1 U1324 ( .A(n744), .B(n1655), .S0(n1656), .Y(\U2/temp_y[2] ) );
  MXI2X1 U1326 ( .A(n745), .B(n2565), .S0(n1660), .Y(\U2/temp_y[1] ) );
  AOI22X1 U1735 ( .A0(temp1t[6]), .A1(temp4t[6]), .B0(n1042), .B1(n1033), .Y(
        n1806) );
  INVX8 U433 ( .A(n1370), .Y(n991) );
  INVX1 U186 ( .A(n2565), .Y(n745) );
  MXI2X1 U943 ( .A(n1354), .B(n992), .S0(n1363), .Y(\U5/Xt[5] ) );
  AOI2BB2X1 U1362 ( .B0(n2557), .B1(n1700), .A0N(n2557), .A1N(n1700), .Y(n1699) );
  MXI2X1 U1092 ( .A(n1464), .B(n965), .S0(n1478), .Y(\U4/Xt[3] ) );
  MXI2X1 U1367 ( .A(n1707), .B(n749), .S0(n1708), .Y(\U2/temp_x[1] ) );
  ADDFX2 \intadd_45/U2  ( .A(\intadd_45/A[8] ), .B(\intadd_39/B[7] ), .CI(
        \intadd_45/n2 ), .CO(\intadd_45/n1 ), .S(\intadd_35/B[5] ) );
  ADDFX2 \intadd_39/U2  ( .A(n2057), .B(\intadd_39/B[8] ), .CI(\intadd_39/n2 ), 
        .CO(\intadd_39/n1 ), .S(\intadd_33/A[5] ) );
  INVX4 U529 ( .A(temp3t[3]), .Y(n1083) );
  CLKINVX3 U486 ( .A(temp4t[5]), .Y(n1041) );
  ADDFX2 \intadd_47/U6  ( .A(n1100), .B(\U5/temp1[4] ), .CI(\intadd_47/n6 ), 
        .CO(\intadd_47/n5 ), .S(\intadd_38/B[3] ) );
  ADDFX2 \intadd_48/U6  ( .A(\U5/temp1[3] ), .B(\U5/temp2[4] ), .CI(
        \intadd_48/n6 ), .CO(\intadd_48/n5 ), .S(\intadd_38/A[0] ) );
  ADDFX2 \intadd_42/U5  ( .A(\intadd_38/A[2] ), .B(n802), .CI(\intadd_42/n5 ), 
        .CO(\intadd_42/n4 ), .S(\U5/temp7[6] ) );
  ADDFX2 \intadd_35/U11  ( .A(\intadd_35/A[0] ), .B(\intadd_35/B[0] ), .CI(
        \intadd_35/CI ), .CO(\intadd_35/n10 ), .S(\intadd_35/SUM[0] ) );
  AOI222X4 U714 ( .A0(x1[1]), .A1(x6[1]), .B0(x1[1]), .B1(n587), .C0(x6[1]), 
        .C1(n587), .Y(n1215) );
  OAI222X4 U705 ( .A0(x1[4]), .A1(x6[4]), .B0(x1[4]), .B1(n583), .C0(x6[4]), 
        .C1(n583), .Y(n1212) );
  AOI222X4 U702 ( .A0(x6[5]), .A1(x1[5]), .B0(x6[5]), .B1(n582), .C0(x1[5]), 
        .C1(n582), .Y(n1211) );
  ADDFX2 \intadd_46/U6  ( .A(\U4/temp1[4] ), .B(\U4/temp2[3] ), .CI(
        \intadd_46/n6 ), .CO(\intadd_46/n5 ), .S(\intadd_37/B[3] ) );
  ADDFX2 \intadd_50/U6  ( .A(n1061), .B(\U4/temp2[3] ), .CI(\intadd_50/n6 ), 
        .CO(\intadd_50/n5 ), .S(\intadd_41/A[2] ) );
  ADDFX2 \intadd_50/U4  ( .A(n1018), .B(\U4/temp2[5] ), .CI(\intadd_50/n4 ), 
        .CO(\intadd_50/n3 ), .S(\intadd_41/A[4] ) );
  AOI222X4 U658 ( .A0(x3[1]), .A1(x4[1]), .B0(x3[1]), .B1(n615), .C0(x4[1]), 
        .C1(n615), .Y(n1197) );
  OAI222X4 U655 ( .A0(x3[2]), .A1(x4[2]), .B0(x3[2]), .B1(n614), .C0(x4[2]), 
        .C1(n614), .Y(n1196) );
  AOI222X4 U652 ( .A0(x4[3]), .A1(x3[3]), .B0(x4[3]), .B1(n613), .C0(x3[3]), 
        .C1(n613), .Y(n1195) );
  AOI222X4 U646 ( .A0(x4[5]), .A1(x3[5]), .B0(x4[5]), .B1(n610), .C0(x3[5]), 
        .C1(n610), .Y(n1193) );
  OAI222X4 U600 ( .A0(n584), .A1(x6[2]), .B0(n584), .B1(n1154), .C0(x6[2]), 
        .C1(n1154), .Y(n1152) );
  OAI222X4 U632 ( .A0(n612), .A1(x4[2]), .B0(n612), .B1(n1186), .C0(x4[2]), 
        .C1(n1186), .Y(n1184) );
  ADDFX2 \intadd_38/U5  ( .A(\intadd_38/A[5] ), .B(\intadd_38/B[5] ), .CI(
        \intadd_38/n5 ), .CO(\intadd_38/n4 ), .S(\intadd_38/SUM[5] ) );
  AND2X2 U836 ( .A(\U1/result6[0] ), .B(\U1/temp_yyyt[0] ), .Y(\intadd_26/CI )
         );
  OAI222X4 U612 ( .A0(n595), .A1(x5[4]), .B0(n595), .B1(n1166), .C0(x5[4]), 
        .C1(n1166), .Y(n1164) );
  OAI222X4 U580 ( .A0(n567), .A1(x7[4]), .B0(n567), .B1(n1134), .C0(x7[4]), 
        .C1(n1134), .Y(n1132) );
  DFFHQX4 \U9/temp_reg[1]  ( .D(temp3[1]), .CK(clk), .Q(temp3t[1]) );
  DFFHQX2 \U8/temp_reg[3]  ( .D(temp2[3]), .CK(clk), .Q(temp2t[3]) );
  DFFHQX4 \U10/temp_reg[6]  ( .D(temp4[6]), .CK(clk), .Q(temp4t[6]) );
  DFFHQX2 \U8/temp_reg[5]  ( .D(temp2[5]), .CK(clk), .Q(temp2t[5]) );
  DFFHQX2 \U3/U20/temp_reg[11]  ( .D(\U3/temp9[11] ), .CK(clk), .Q(
        \U3/temp12[1] ) );
  DFFHQX2 \U3/U21/temp_reg[10]  ( .D(n680), .CK(clk), .Q(\U3/temp11[0] ) );
  DFFHQX2 \U13/temp_reg[9]  ( .D(temp7[9]), .CK(clk), .Q(\U4/temp2[9] ) );
  DFFHQX2 \U11/temp_reg[5]  ( .D(temp5[5]), .CK(clk), .Q(\U5/temp1[4] ) );
  DFFHQX2 \U11/temp_reg[3]  ( .D(temp5[3]), .CK(clk), .Q(\U5/temp1[2] ) );
  DFFHQX2 \U4/U11/temp_reg[9]  ( .D(\U4/temp5[9] ), .CK(clk), .Q(
        \U4/U5/temp[6] ) );
  DFFHQX2 \U5/U12/temp_reg[9]  ( .D(\U5/temp7[9] ), .CK(clk), .Q(
        \U5/U6/temp[6] ) );
  DFFHQX2 \U5/U11/temp_reg[9]  ( .D(n789), .CK(clk), .Q(\U5/U5/temp[6] ) );
  DFFHQX2 \U4/U12/temp_reg[9]  ( .D(n813), .CK(clk), .Q(\U4/U6/temp[6] ) );
  DFFHQX2 \U11/temp_reg[7]  ( .D(temp5[7]), .CK(clk), .Q(\U5/temp1[6] ) );
  DFFHQX2 \U14/temp_reg[9]  ( .D(temp8[9]), .CK(clk), .Q(\U5/temp2[9] ) );
  DFFHQX2 \U5/U12/temp_reg[7]  ( .D(\U5/temp7[7] ), .CK(clk), .Q(
        \U5/U6/temp[4] ) );
  DFFHQX2 \U5/U11/temp_reg[7]  ( .D(n791), .CK(clk), .Q(\U5/U5/temp[4] ) );
  DFFHQX2 \U4/U12/temp_reg[7]  ( .D(n815), .CK(clk), .Q(\U4/U6/temp[4] ) );
  DFFHQX2 \U4/U11/temp_reg[7]  ( .D(\U4/temp5[7] ), .CK(clk), .Q(
        \U4/U5/temp[4] ) );
  DFFHQX1 \U2/U20/temp_reg[10]  ( .D(\U2/temp_x[10] ), .CK(clk), .Q(
        \U2/result1[9] ) );
  DFFHQX2 \U7/temp_reg[5]  ( .D(temp1[5]), .CK(clk), .Q(temp1t[5]) );
  DFFHQX2 \U3/U21/temp_reg[3]  ( .D(n708), .CK(clk), .Q(\U3/temp10t[3] ) );
  DFFHQX2 \U3/U21/temp_reg[2]  ( .D(n712), .CK(clk), .Q(\U3/temp10t[2] ) );
  DFFHQX2 \U9/temp_reg[4]  ( .D(temp3[4]), .CK(clk), .Q(temp3t[4]) );
  DFFHQX2 \U14/temp_reg[2]  ( .D(temp8[2]), .CK(clk), .Q(\U5/temp2[1] ) );
  DFFHQX2 \U3/U21/temp_reg[5]  ( .D(n700), .CK(clk), .Q(\U3/temp10t[5] ) );
  DFFHQX2 \U3/U21/temp_reg[9]  ( .D(n685), .CK(clk), .Q(\U3/temp10t[9] ) );
  DFFHQX2 \U3/U21/temp_reg[7]  ( .D(n687), .CK(clk), .Q(\U3/temp10t[7] ) );
  DFFHQX2 \U7/temp_reg[7]  ( .D(temp1[7]), .CK(clk), .Q(temp1t[7]) );
  DFFHQX2 \U9/temp_reg[8]  ( .D(temp3[8]), .CK(clk), .Q(temp3t[8]) );
  DFFHQX2 \U7/temp_reg[9]  ( .D(temp1[9]), .CK(clk), .Q(temp1t[9]) );
  DFFHQX2 \U9/temp_reg[9]  ( .D(temp3[9]), .CK(clk), .Q(temp3t[9]) );
  DFFHQX2 \U10/temp_reg[8]  ( .D(temp4[8]), .CK(clk), .Q(temp4t[8]) );
  DFFHQX1 \U2/U21/temp_reg[10]  ( .D(\U2/temp_y[10] ), .CK(clk), .Q(
        \U2/result2[9] ) );
  DFFHQX2 \U6/U8/temp_reg[10]  ( .D(\intadd_40/n1 ), .CK(clk), .Q(
        \U6/temp6[10] ) );
  DFFHQX2 \U3/U21/temp_reg[8]  ( .D(n686), .CK(clk), .Q(\U3/temp10t[8] ) );
  DFFHQX2 \U14/temp_reg[3]  ( .D(temp8[3]), .CK(clk), .Q(\U5/temp2[2] ) );
  DFFHQX2 \U5/U11/temp_reg[11]  ( .D(\U5/temp5[11] ), .CK(clk), .Q(
        \U5/U5/temp[11] ) );
  DFFHQX2 \U5/U12/temp_reg[11]  ( .D(\U5/temp7[11] ), .CK(clk), .Q(
        \U5/U6/temp[11] ) );
  DFFHQX2 \U4/U12/temp_reg[11]  ( .D(\U4/temp7[11] ), .CK(clk), .Q(
        \U4/U6/temp[11] ) );
  DFFHQX2 \U4/U11/temp_reg[11]  ( .D(\U4/temp5[11] ), .CK(clk), .Q(
        \U4/U5/temp[11] ) );
  DFFHQX2 \U14/temp_reg[5]  ( .D(temp8[5]), .CK(clk), .Q(\U5/temp2[4] ) );
  DFFHQX2 \U3/U21/temp_reg[4]  ( .D(n704), .CK(clk), .Q(\U3/temp10t[4] ) );
  DFFHQX2 \U3/U21/temp_reg[6]  ( .D(n696), .CK(clk), .Q(\U3/temp10t[6] ) );
  CLKINVX3 U501 ( .A(\U5/temp1[7] ), .Y(n1056) );
  CLKINVX3 U540 ( .A(\U5/temp1[5] ), .Y(n1094) );
  ADDFX2 \intadd_36/U11  ( .A(n921), .B(\U6/temp5[1] ), .CI(\intadd_36/CI ), 
        .CO(\intadd_36/n10 ), .S(\intadd_36/SUM[0] ) );
  AOI2BB2X2 U820 ( .B0(\U5/temp2[9] ), .B1(n1117), .A0N(n1117), .A1N(
        \U5/temp2[9] ), .Y(n1244) );
  ADDFX2 \intadd_25/U21  ( .A(\U1/result5[1] ), .B(\U1/temp_xxxt[1] ), .CI(
        \intadd_25/CI ), .CO(\intadd_25/n20 ), .S(\intadd_25/SUM[0] ) );
  ADDFX2 \intadd_26/U21  ( .A(\U1/result6[1] ), .B(\U1/temp_yyyt[1] ), .CI(
        \intadd_26/CI ), .CO(\intadd_26/n20 ), .S(\intadd_26/SUM[0] ) );
  ADDFX2 \intadd_40/U10  ( .A(n1055), .B(\U4/temp1[3] ), .CI(\intadd_40/CI ), 
        .CO(\intadd_40/n9 ), .S(\intadd_40/SUM[0] ) );
  ADDFX2 \intadd_29/U12  ( .A(result3[1]), .B(result1[1]), .CI(\intadd_29/CI ), 
        .CO(\intadd_29/n11 ), .S(s4[1]) );
  ADDFX2 \intadd_26/U20  ( .A(\U1/result6[2] ), .B(\U1/temp_yyyt[2] ), .CI(
        \intadd_26/n20 ), .CO(\intadd_26/n19 ), .S(\intadd_26/SUM[1] ) );
  ADDFX2 \intadd_25/U20  ( .A(\U1/result5[2] ), .B(\U1/temp_xxxt[2] ), .CI(
        \intadd_25/n20 ), .CO(\intadd_25/n19 ), .S(\intadd_25/SUM[1] ) );
  ADDFX2 \intadd_48/U9  ( .A(\U5/temp1[0] ), .B(\U5/temp2[1] ), .CI(
        \intadd_48/CI ), .CO(\intadd_48/n8 ), .S(\intadd_42/B[0] ) );
  ADDFX2 \intadd_50/U8  ( .A(n1110), .B(\U4/temp2[1] ), .CI(\intadd_50/CI ), 
        .CO(\intadd_50/n7 ), .S(\intadd_41/A[0] ) );
  ADDFX2 \intadd_47/U9  ( .A(n852), .B(\U5/temp1[1] ), .CI(\intadd_47/CI ), 
        .CO(\intadd_47/n8 ), .S(\intadd_38/CI ) );
  ADDFX2 \intadd_34/U11  ( .A(\U6/temp6[1] ), .B(\U6/temp3t[1] ), .CI(
        \intadd_34/CI ), .CO(\intadd_34/n10 ), .S(\U6/Xt[0] ) );
  ADDFX2 \intadd_36/U10  ( .A(n906), .B(\U6/temp5[2] ), .CI(\intadd_36/n10 ), 
        .CO(\intadd_36/n9 ), .S(\intadd_36/SUM[1] ) );
  ADDFX2 \intadd_30/U12  ( .A(result4[1]), .B(result2[1]), .CI(\intadd_30/CI ), 
        .CO(\intadd_30/n11 ), .S(s5[1]) );
  ADDFX2 \intadd_44/U10  ( .A(n2068), .B(\intadd_44/B[0] ), .CI(\intadd_44/CI ), .CO(\intadd_44/n9 ), .S(\U2/Ytt[0] ) );
  ADDFX2 \intadd_49/U8  ( .A(\U4/temp1[0] ), .B(\U4/temp2[3] ), .CI(
        \intadd_49/CI ), .CO(\intadd_49/n7 ), .S(\U6/temp3[1] ) );
  ADDFX2 \intadd_40/U9  ( .A(n1057), .B(\U4/temp1[4] ), .CI(\intadd_40/n9 ), 
        .CO(\intadd_40/n8 ), .S(\intadd_40/SUM[1] ) );
  ADDFX2 \intadd_43/U10  ( .A(n2067), .B(\intadd_43/B[0] ), .CI(\intadd_43/CI ), .CO(\intadd_43/n9 ), .S(\U2/Xtt[0] ) );
  ADDFX2 \intadd_29/U11  ( .A(result3[2]), .B(result1[2]), .CI(\intadd_29/n11 ), .CO(\intadd_29/n10 ), .S(s4[2]) );
  ADDFX2 \intadd_36/U9  ( .A(n907), .B(\U6/temp5[3] ), .CI(\intadd_36/n9 ), 
        .CO(\intadd_36/n8 ), .S(\intadd_36/SUM[2] ) );
  ADDFX2 \intadd_46/U9  ( .A(\U4/temp1[1] ), .B(\U4/temp2[0] ), .CI(
        \intadd_46/CI ), .CO(\intadd_46/n8 ), .S(\intadd_37/CI ) );
  ADDFX2 \intadd_50/U7  ( .A(n1059), .B(\U4/temp2[2] ), .CI(\intadd_50/n7 ), 
        .CO(\intadd_50/n6 ), .S(\intadd_41/A[1] ) );
  ADDFX2 \intadd_48/U8  ( .A(\U5/temp1[1] ), .B(\U5/temp2[2] ), .CI(
        \intadd_48/n8 ), .CO(\intadd_48/n7 ), .S(\intadd_42/A[1] ) );
  ADDFX2 \intadd_31/U11  ( .A(result7[1]), .B(n915), .CI(n927), .CO(
        \intadd_31/n10 ), .S(\intadd_31/SUM[0] ) );
  ADDFX2 \intadd_30/U11  ( .A(result4[2]), .B(result2[2]), .CI(\intadd_30/n11 ), .CO(\intadd_30/n10 ), .S(s5[2]) );
  ADDFX2 \intadd_47/U8  ( .A(n1099), .B(\U5/temp1[2] ), .CI(\intadd_47/n8 ), 
        .CO(\intadd_47/n7 ), .S(\intadd_38/B[1] ) );
  ADDFX2 \intadd_26/U19  ( .A(\U1/result6[13] ), .B(\U1/temp_yyyt[3] ), .CI(
        \intadd_26/n19 ), .CO(\intadd_26/n18 ), .S(\intadd_26/SUM[2] ) );
  ADDFX2 \intadd_32/U11  ( .A(result8[1]), .B(n918), .CI(n928), .CO(
        \intadd_32/n10 ), .S(\intadd_32/SUM[0] ) );
  ADDFX2 \intadd_34/U10  ( .A(\U6/temp6[2] ), .B(\U6/temp3t[2] ), .CI(
        \intadd_34/n10 ), .CO(\intadd_34/n9 ), .S(\U6/Xt[1] ) );
  ADDFX2 \intadd_25/U19  ( .A(\U1/result5[13] ), .B(\U1/temp_xxxt[3] ), .CI(
        \intadd_25/n19 ), .CO(\intadd_25/n18 ), .S(\intadd_25/SUM[2] ) );
  INVX2 U12 ( .A(n1223), .Y(n571) );
  ADDFX2 \intadd_34/U9  ( .A(\U6/temp6[3] ), .B(\U6/temp3t[3] ), .CI(
        \intadd_34/n9 ), .CO(\intadd_34/n8 ), .S(\U6/Xt[2] ) );
  ADDFX2 \intadd_36/U8  ( .A(\U6/temp5[4] ), .B(n926), .CI(\intadd_36/n8 ), 
        .CO(\intadd_36/n7 ), .S(\intadd_36/SUM[3] ) );
  ADDFX2 \intadd_46/U8  ( .A(\U4/temp1[2] ), .B(\U4/temp2[1] ), .CI(
        \intadd_46/n8 ), .CO(\intadd_46/n7 ), .S(\intadd_37/B[1] ) );
  ADDFX2 \intadd_32/U10  ( .A(result8[2]), .B(n919), .CI(\intadd_32/n10 ), 
        .CO(\intadd_32/n9 ), .S(\intadd_32/SUM[1] ) );
  ADDFX2 \intadd_40/U8  ( .A(n1058), .B(\U4/temp1[5] ), .CI(\intadd_40/n8 ), 
        .CO(\intadd_40/n7 ), .S(\intadd_40/SUM[2] ) );
  ADDFX2 \intadd_26/U18  ( .A(\U1/result6[13] ), .B(\U1/temp_yyyt[4] ), .CI(
        \intadd_26/n18 ), .CO(\intadd_26/n17 ), .S(\intadd_26/SUM[3] ) );
  ADDFX2 \intadd_49/U7  ( .A(\U4/temp1[1] ), .B(\U4/temp2[4] ), .CI(
        \intadd_49/n7 ), .CO(\intadd_49/n6 ), .S(\U6/temp3[2] ) );
  ADDFX2 \intadd_30/U10  ( .A(result4[3]), .B(result2[3]), .CI(\intadd_30/n10 ), .CO(\intadd_30/n9 ), .S(s5[3]) );
  ADDFX2 \intadd_29/U10  ( .A(result3[3]), .B(result1[3]), .CI(\intadd_29/n10 ), .CO(\intadd_29/n9 ), .S(s4[3]) );
  ADDFX2 \intadd_31/U10  ( .A(result7[2]), .B(n916), .CI(\intadd_31/n10 ), 
        .CO(\intadd_31/n9 ), .S(\intadd_31/SUM[1] ) );
  ADDFX2 \intadd_25/U18  ( .A(\U1/result5[13] ), .B(\U1/temp_xxxt[4] ), .CI(
        \intadd_25/n18 ), .CO(\intadd_25/n17 ), .S(\intadd_25/SUM[3] ) );
  AOI222X4 U680 ( .A0(x5[3]), .A1(x2[3]), .B0(x5[3]), .B1(n599), .C0(x2[3]), 
        .C1(n599), .Y(n1204) );
  ADDFX2 \intadd_30/U9  ( .A(result4[4]), .B(result2[4]), .CI(\intadd_30/n9 ), 
        .CO(\intadd_30/n8 ), .S(s5[4]) );
  ADDFX2 \intadd_32/U9  ( .A(result8[3]), .B(n900), .CI(\intadd_32/n9 ), .CO(
        \intadd_32/n8 ), .S(\intadd_32/SUM[2] ) );
  ADDFX2 \intadd_26/U17  ( .A(\U1/temp_yyyt[5] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n17 ), .CO(\intadd_26/n16 ), .S(\intadd_26/SUM[4] ) );
  ADDFX2 \intadd_43/U9  ( .A(\intadd_43/A[1] ), .B(\intadd_43/B[1] ), .CI(
        \intadd_43/n9 ), .CO(\intadd_43/n8 ), .S(\U2/Xtt[1] ) );
  ADDFX2 \intadd_40/U7  ( .A(n1014), .B(\U4/temp1[6] ), .CI(\intadd_40/n7 ), 
        .CO(\intadd_40/n6 ), .S(\intadd_40/SUM[3] ) );
  ADDFX2 \intadd_34/U8  ( .A(\U6/temp6[4] ), .B(\U6/temp5[0] ), .CI(
        \intadd_34/n8 ), .CO(\intadd_34/n7 ), .S(\U6/Xt[3] ) );
  ADDFX2 \intadd_36/U7  ( .A(\U6/temp5[5] ), .B(n929), .CI(\intadd_36/n7 ), 
        .CO(\intadd_36/n6 ), .S(\intadd_36/SUM[4] ) );
  NOR2X4 U1548 ( .A(n930), .B(n1258), .Y(n1234) );
  ADDFX2 \intadd_29/U9  ( .A(result3[4]), .B(result1[4]), .CI(\intadd_29/n9 ), 
        .CO(\intadd_29/n8 ), .S(s4[4]) );
  ADDFX2 \intadd_49/U6  ( .A(\U4/temp1[2] ), .B(\U4/temp2[5] ), .CI(
        \intadd_49/n6 ), .CO(\intadd_49/n5 ), .S(\U6/temp3[3] ) );
  ADDFX2 \intadd_31/U9  ( .A(result7[3]), .B(n895), .CI(\intadd_31/n9 ), .CO(
        \intadd_31/n8 ), .S(\intadd_31/SUM[2] ) );
  ADDFX2 \intadd_50/U5  ( .A(n1017), .B(\U4/temp2[4] ), .CI(\intadd_50/n5 ), 
        .CO(\intadd_50/n4 ), .S(\intadd_41/A[3] ) );
  ADDFX2 \intadd_44/U9  ( .A(\intadd_44/A[1] ), .B(\intadd_44/B[1] ), .CI(
        \intadd_44/n9 ), .CO(\intadd_44/n8 ), .S(\U2/Ytt[1] ) );
  NOR2X4 U1537 ( .A(n931), .B(n1252), .Y(n1233) );
  ADDFX2 \intadd_25/U17  ( .A(\U1/temp_xxxt[5] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n17 ), .CO(\intadd_25/n16 ), .S(\intadd_25/SUM[4] ) );
  ADDFX2 \intadd_26/U16  ( .A(\U1/temp_yyyt[6] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n16 ), .CO(\intadd_26/n15 ), .S(\intadd_26/SUM[5] ) );
  ADDFX2 \intadd_34/U7  ( .A(\U6/temp6[5] ), .B(\U6/temp5[1] ), .CI(
        \intadd_34/n7 ), .CO(\intadd_34/n6 ), .S(\U6/Xt[4] ) );
  ADDFX2 \intadd_36/U6  ( .A(n885), .B(\U6/temp6[2] ), .CI(\intadd_36/n6 ), 
        .CO(\intadd_36/n5 ), .S(\intadd_36/SUM[5] ) );
  ADDFX2 \intadd_32/U8  ( .A(result8[4]), .B(n901), .CI(\intadd_32/n8 ), .CO(
        \intadd_32/n7 ), .S(\intadd_32/SUM[3] ) );
  ADDFX2 \intadd_43/U8  ( .A(n2067), .B(n2066), .CI(\intadd_43/n8 ), .CO(
        \intadd_43/n7 ), .S(\U2/Xtt[2] ) );
  ADDFX2 \intadd_44/U8  ( .A(n2068), .B(n2065), .CI(\intadd_44/n8 ), .CO(
        \intadd_44/n7 ), .S(\U2/Ytt[2] ) );
  ADDFX2 \intadd_29/U8  ( .A(result3[5]), .B(result1[5]), .CI(\intadd_29/n8 ), 
        .CO(\intadd_29/n7 ), .S(s4[5]) );
  ADDFX2 \intadd_49/U5  ( .A(\U4/temp1[3] ), .B(\U4/temp2[6] ), .CI(
        \intadd_49/n5 ), .CO(\intadd_49/n4 ), .S(\U6/temp3[4] ) );
  ADDFX2 \intadd_40/U6  ( .A(n1015), .B(\U4/temp1[7] ), .CI(\intadd_40/n6 ), 
        .CO(\intadd_40/n5 ), .S(\intadd_40/SUM[4] ) );
  ADDFX2 \intadd_25/U16  ( .A(\U1/temp_xxxt[6] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n16 ), .CO(\intadd_25/n15 ), .S(\intadd_25/SUM[5] ) );
  ADDFX2 \intadd_31/U8  ( .A(result7[4]), .B(n896), .CI(\intadd_31/n8 ), .CO(
        \intadd_31/n7 ), .S(\intadd_31/SUM[3] ) );
  ADDFX2 \intadd_30/U8  ( .A(result4[5]), .B(result2[5]), .CI(\intadd_30/n8 ), 
        .CO(\intadd_30/n7 ), .S(s5[5]) );
  ADDFX2 \intadd_29/U7  ( .A(result3[6]), .B(result1[6]), .CI(\intadd_29/n7 ), 
        .CO(\intadd_29/n6 ), .S(s4[6]) );
  ADDFX2 \intadd_34/U6  ( .A(\U6/temp5[2] ), .B(\U6/temp6[10] ), .CI(
        \intadd_34/n6 ), .CO(\intadd_34/n5 ), .S(\U6/Xt[5] ) );
  ADDFX2 \intadd_44/U7  ( .A(\intadd_44/B[1] ), .B(\intadd_44/B[3] ), .CI(
        \intadd_44/n7 ), .CO(\intadd_44/n6 ), .S(\U2/Ytt[3] ) );
  ADDFX2 \intadd_37/U10  ( .A(n829), .B(\intadd_37/B[0] ), .CI(\intadd_37/CI ), 
        .CO(\intadd_37/n9 ), .S(\U4/temp5[1] ) );
  ADDFX2 \intadd_38/U10  ( .A(\intadd_38/A[0] ), .B(\intadd_38/B[0] ), .CI(
        \intadd_38/CI ), .CO(\intadd_38/n9 ), .S(\intadd_38/SUM[0] ) );
  ADDFX2 \intadd_40/U5  ( .A(\U4/temp2[5] ), .B(n1119), .CI(\intadd_40/n5 ), 
        .CO(\intadd_40/n4 ), .S(\intadd_40/SUM[5] ) );
  ADDFX2 \intadd_36/U5  ( .A(n910), .B(\U6/temp6[3] ), .CI(\intadd_36/n5 ), 
        .CO(\intadd_36/n4 ), .S(\intadd_36/SUM[6] ) );
  ADDFX2 \intadd_49/U4  ( .A(\U4/temp1[4] ), .B(\U4/temp2[7] ), .CI(
        \intadd_49/n4 ), .CO(\intadd_49/n3 ), .S(\U6/temp3[5] ) );
  ADDFX2 \intadd_43/U7  ( .A(\intadd_43/B[1] ), .B(\intadd_43/B[3] ), .CI(
        \intadd_43/n7 ), .CO(\intadd_43/n6 ), .S(\U2/Xtt[3] ) );
  ADDFX2 \intadd_45/U10  ( .A(n786), .B(\intadd_45/B[0] ), .CI(\intadd_45/CI ), 
        .CO(\intadd_45/n9 ), .S(\intadd_45/SUM[0] ) );
  ADDFX2 \intadd_25/U15  ( .A(\U1/temp_xxxt[7] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n15 ), .CO(\intadd_25/n14 ), .S(\intadd_25/SUM[6] ) );
  ADDFX2 \intadd_42/U10  ( .A(\intadd_42/A[0] ), .B(\intadd_42/B[0] ), .CI(
        n809), .CO(\intadd_42/n9 ), .S(\U5/temp7[1] ) );
  ADDFX2 \intadd_32/U7  ( .A(result8[5]), .B(n902), .CI(\intadd_32/n7 ), .CO(
        \intadd_32/n6 ), .S(\intadd_32/SUM[4] ) );
  ADDFX2 \intadd_31/U7  ( .A(result7[5]), .B(n897), .CI(\intadd_31/n7 ), .CO(
        \intadd_31/n6 ), .S(\intadd_31/SUM[4] ) );
  ADDFX2 \intadd_30/U7  ( .A(result4[6]), .B(result2[6]), .CI(\intadd_30/n7 ), 
        .CO(\intadd_30/n6 ), .S(s5[6]) );
  ADDFX2 \intadd_26/U15  ( .A(\U1/temp_yyyt[7] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n15 ), .CO(\intadd_26/n14 ), .S(\intadd_26/SUM[6] ) );
  ADDFX2 \intadd_31/U6  ( .A(result7[6]), .B(n871), .CI(\intadd_31/n6 ), .CO(
        \intadd_31/n5 ), .S(\intadd_31/SUM[5] ) );
  ADDFX2 \intadd_43/U6  ( .A(n2066), .B(n2064), .CI(\intadd_43/n6 ), .CO(
        \intadd_43/n5 ), .S(\U2/Xtt[4] ) );
  ADDFX2 \intadd_40/U4  ( .A(n1024), .B(\U4/temp2[6] ), .CI(\intadd_40/n4 ), 
        .CO(\intadd_40/n3 ), .S(\intadd_40/SUM[6] ) );
  ADDFX2 \intadd_49/U3  ( .A(\U4/temp2[9] ), .B(\U4/temp1[5] ), .CI(
        \intadd_49/n3 ), .CO(\intadd_49/n2 ), .S(\U6/temp3[6] ) );
  ADDFX2 \intadd_39/U10  ( .A(\intadd_39/A[0] ), .B(n2050), .CI(\intadd_39/CI ), .CO(\intadd_39/n9 ), .S(\intadd_35/A[0] ) );
  ADDFX2 \intadd_30/U6  ( .A(result4[7]), .B(result2[7]), .CI(\intadd_30/n6 ), 
        .CO(\intadd_30/n5 ), .S(s5[7]) );
  ADDFX2 \intadd_42/U9  ( .A(\intadd_42/A[1] ), .B(n808), .CI(\intadd_42/n9 ), 
        .CO(\intadd_42/n8 ), .S(\U5/temp7[2] ) );
  ADDFX2 U479 ( .A(n2065), .B(n2063), .CI(\intadd_44/n6 ), .CO(\intadd_44/n5 ), 
        .S(\U2/Ytt[4] ) );
  ADDFX2 \intadd_32/U6  ( .A(result8[6]), .B(n876), .CI(\intadd_32/n6 ), .CO(
        \intadd_32/n5 ), .S(\intadd_32/SUM[5] ) );
  ADDFX2 \intadd_34/U5  ( .A(\U6/temp5[3] ), .B(\U6/temp6[10] ), .CI(
        \intadd_34/n5 ), .CO(\intadd_34/n4 ), .S(\U6/Xt[6] ) );
  ADDFX2 \intadd_26/U14  ( .A(\U1/result6[0] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n14 ), .CO(\intadd_26/n13 ), .S(\intadd_26/SUM[7] ) );
  ADDFX2 \intadd_29/U6  ( .A(result3[7]), .B(result1[7]), .CI(\intadd_29/n6 ), 
        .CO(\intadd_29/n5 ), .S(s4[7]) );
  ADDFX2 \intadd_37/U9  ( .A(n828), .B(\intadd_37/B[1] ), .CI(\intadd_37/n9 ), 
        .CO(\intadd_37/n8 ), .S(\U4/temp5[2] ) );
  ADDFX2 \intadd_41/U10  ( .A(\intadd_41/A[0] ), .B(\intadd_41/B[0] ), .CI(
        \intadd_37/B[3] ), .CO(\intadd_41/n9 ), .S(\intadd_41/SUM[0] ) );
  ADDFX2 \intadd_38/U9  ( .A(\intadd_38/A[1] ), .B(\intadd_38/B[1] ), .CI(
        \intadd_38/n9 ), .CO(\intadd_38/n8 ), .S(\intadd_38/SUM[1] ) );
  ADDFX2 \intadd_36/U4  ( .A(n911), .B(\U6/temp6[4] ), .CI(\intadd_36/n4 ), 
        .CO(\intadd_36/n3 ), .S(\intadd_36/SUM[7] ) );
  ADDFX2 \intadd_37/U8  ( .A(n827), .B(\intadd_37/B[2] ), .CI(\intadd_37/n8 ), 
        .CO(\intadd_37/n7 ), .S(\U4/temp5[3] ) );
  ADDFX2 \intadd_49/U2  ( .A(\U4/temp2[9] ), .B(\U4/temp1[6] ), .CI(
        \intadd_49/n2 ), .CO(\intadd_49/n1 ), .S(\U6/temp3[7] ) );
  ADDFX2 \intadd_41/U9  ( .A(\intadd_41/A[1] ), .B(\intadd_37/B[4] ), .CI(
        \intadd_41/n9 ), .CO(\intadd_41/n8 ), .S(\intadd_41/SUM[1] ) );
  ADDFX2 \intadd_40/U3  ( .A(n1023), .B(\U4/temp2[7] ), .CI(\intadd_40/n3 ), 
        .CO(\intadd_40/n2 ), .S(\intadd_40/SUM[7] ) );
  ADDFX2 \intadd_42/U8  ( .A(\intadd_42/A[2] ), .B(n807), .CI(\intadd_42/n8 ), 
        .CO(\intadd_42/n7 ), .S(\U5/temp7[3] ) );
  ADDFX2 \intadd_36/U3  ( .A(n912), .B(\U6/temp6[5] ), .CI(\intadd_36/n3 ), 
        .CO(\intadd_36/n2 ), .S(\intadd_36/SUM[8] ) );
  ADDFX2 \intadd_34/U4  ( .A(\U6/temp5[4] ), .B(\U6/temp6[10] ), .CI(
        \intadd_34/n4 ), .CO(\intadd_34/n3 ), .S(\U6/Xt[7] ) );
  ADDFX2 \intadd_43/U5  ( .A(\intadd_43/B[3] ), .B(\intadd_43/B[5] ), .CI(
        \intadd_43/n5 ), .CO(\intadd_43/n4 ), .S(\U2/Xtt[5] ) );
  ADDFX2 \intadd_44/U5  ( .A(\intadd_44/B[3] ), .B(n2158), .CI(\intadd_44/n5 ), 
        .CO(\intadd_44/n4 ), .S(\U2/Ytt[5] ) );
  ADDFX2 \intadd_38/U8  ( .A(\intadd_38/A[2] ), .B(\intadd_38/B[2] ), .CI(
        \intadd_38/n8 ), .CO(\intadd_38/n7 ), .S(\intadd_38/SUM[2] ) );
  ADDFX2 \intadd_32/U5  ( .A(result8[7]), .B(n877), .CI(\intadd_32/n5 ), .CO(
        \intadd_32/n4 ), .S(\intadd_32/SUM[6] ) );
  ADDFX2 \intadd_30/U5  ( .A(result4[8]), .B(result2[8]), .CI(\intadd_30/n5 ), 
        .CO(\intadd_30/n4 ), .S(s5[8]) );
  ADDFX2 \intadd_29/U5  ( .A(result3[8]), .B(result1[8]), .CI(\intadd_29/n5 ), 
        .CO(\intadd_29/n4 ), .S(s4[8]) );
  ADDFX2 \intadd_39/U9  ( .A(\intadd_39/A[1] ), .B(\intadd_39/B[1] ), .CI(
        \intadd_39/n9 ), .CO(\intadd_39/n8 ), .S(\intadd_35/A[1] ) );
  ADDFX2 \intadd_31/U5  ( .A(result7[7]), .B(n872), .CI(\intadd_31/n5 ), .CO(
        \intadd_31/n4 ), .S(\intadd_31/SUM[6] ) );
  ADDFX2 \intadd_45/U9  ( .A(n784), .B(\intadd_39/CI ), .CI(\intadd_45/n9 ), 
        .CO(\intadd_45/n8 ), .S(\intadd_45/SUM[1] ) );
  ADDFX2 U478 ( .A(n2063), .B(n2061), .CI(\intadd_44/n4 ), .CO(\intadd_44/n3 ), 
        .S(\U2/Ytt[6] ) );
  ADDFX2 \intadd_36/U2  ( .A(\U6/temp6[10] ), .B(n891), .CI(\intadd_36/n2 ), 
        .CO(\intadd_36/n1 ), .S(\intadd_36/SUM[9] ) );
  ADDFX2 \intadd_42/U7  ( .A(\intadd_38/A[0] ), .B(n806), .CI(\intadd_42/n7 ), 
        .CO(\intadd_42/n6 ), .S(\U5/temp7[4] ) );
  ADDFX2 \intadd_34/U3  ( .A(\U6/temp5[5] ), .B(\U6/temp6[10] ), .CI(
        \intadd_34/n3 ), .CO(\intadd_34/n2 ), .S(\U6/Xt[8] ) );
  ADDFX2 \intadd_38/U7  ( .A(\intadd_38/A[3] ), .B(\intadd_38/B[3] ), .CI(
        \intadd_38/n7 ), .CO(\intadd_38/n6 ), .S(\intadd_38/SUM[3] ) );
  ADDFX2 \intadd_37/U7  ( .A(n826), .B(\intadd_37/B[3] ), .CI(\intadd_37/n7 ), 
        .CO(\intadd_37/n6 ), .S(\U4/temp5[4] ) );
  ADDFX2 \intadd_43/U4  ( .A(n2064), .B(n2062), .CI(\intadd_43/n4 ), .CO(
        \intadd_43/n3 ), .S(\U2/Xtt[6] ) );
  ADDFX2 \intadd_40/U2  ( .A(\U4/temp2[9] ), .B(n935), .CI(\intadd_40/n2 ), 
        .CO(\intadd_40/n1 ), .S(\intadd_40/SUM[8] ) );
  ADDFX2 \intadd_41/U8  ( .A(\intadd_41/A[2] ), .B(\intadd_37/B[5] ), .CI(
        \intadd_41/n8 ), .CO(\intadd_41/n7 ), .S(\intadd_41/SUM[2] ) );
  ADDFX2 \intadd_30/U4  ( .A(result4[9]), .B(result2[9]), .CI(\intadd_30/n4 ), 
        .CO(\intadd_30/n3 ), .S(s5[9]) );
  ADDFX2 \intadd_32/U4  ( .A(result8[8]), .B(n878), .CI(\intadd_32/n4 ), .CO(
        \intadd_32/n3 ), .S(\intadd_32/SUM[7] ) );
  ADDFX2 \intadd_31/U4  ( .A(result7[8]), .B(n873), .CI(\intadd_31/n4 ), .CO(
        \intadd_31/n3 ), .S(\intadd_31/SUM[7] ) );
  ADDFX2 \intadd_29/U4  ( .A(result3[9]), .B(result1[9]), .CI(\intadd_29/n4 ), 
        .CO(\intadd_29/n3 ), .S(s4[9]) );
  OAI222X4 U727 ( .A0(x0[6]), .A1(x7[6]), .B0(x0[6]), .B1(n566), .C0(x7[6]), 
        .C1(n566), .Y(n1219) );
  ADDFX2 \intadd_42/U6  ( .A(\intadd_38/A[1] ), .B(n805), .CI(\intadd_42/n6 ), 
        .CO(\intadd_42/n5 ), .S(\U5/temp7[5] ) );
  ADDFX2 \intadd_32/U3  ( .A(result8[9]), .B(n862), .CI(\intadd_32/n3 ), .CO(
        \intadd_32/n2 ), .S(\intadd_32/SUM[8] ) );
  ADDFX2 \intadd_37/U6  ( .A(n824), .B(\intadd_37/B[4] ), .CI(\intadd_37/n6 ), 
        .CO(\intadd_37/n5 ), .S(\U4/temp5[5] ) );
  ADDFX2 \intadd_51/U4  ( .A(\intadd_25/SUM[9] ), .B(\intadd_51/B[0] ), .CI(
        \intadd_25/SUM[0] ), .CO(\intadd_51/n3 ), .S(\U1/Xtt[0] ) );
  ADDFX2 \intadd_38/U6  ( .A(\intadd_38/A[4] ), .B(\intadd_38/B[4] ), .CI(
        \intadd_38/n6 ), .CO(\intadd_38/n5 ), .S(\intadd_38/SUM[4] ) );
  ADDFX2 \intadd_30/U3  ( .A(result4[11]), .B(result2[10]), .CI(\intadd_30/n3 ), .CO(\intadd_30/n2 ), .S(s5[10]) );
  ADDFX2 \intadd_44/U3  ( .A(\intadd_44/A[7] ), .B(n2158), .CI(\intadd_44/n3 ), 
        .CO(\intadd_44/n2 ), .S(\U2/Ytt[7] ) );
  ADDFX2 \intadd_31/U3  ( .A(result7[9]), .B(n859), .CI(\intadd_31/n3 ), .CO(
        \intadd_31/n2 ), .S(\intadd_31/SUM[8] ) );
  ADDFX2 \intadd_29/U3  ( .A(result3[11]), .B(result1[10]), .CI(\intadd_29/n3 ), .CO(\intadd_29/n2 ), .S(s4[10]) );
  ADDFX2 \intadd_34/U2  ( .A(n1120), .B(n885), .CI(\intadd_34/n2 ), .CO(
        \intadd_34/n1 ), .S(\U6/Xt[9] ) );
  ADDFX2 \intadd_41/U7  ( .A(\intadd_41/A[3] ), .B(\intadd_37/B[6] ), .CI(
        \intadd_41/n7 ), .CO(\intadd_41/n6 ), .S(\intadd_41/SUM[3] ) );
  ADDFX2 \intadd_43/U3  ( .A(\intadd_43/A[7] ), .B(\intadd_43/B[5] ), .CI(
        \intadd_43/n3 ), .CO(\intadd_43/n2 ), .S(\U2/Xtt[7] ) );
  ADDFX2 \intadd_31/U2  ( .A(result5[11]), .B(n863), .CI(\intadd_31/n2 ), .CO(
        \intadd_31/n1 ), .S(\intadd_31/SUM[9] ) );
  ADDFX2 \intadd_29/U2  ( .A(n854), .B(n867), .CI(\intadd_29/n2 ), .CO(
        \intadd_29/n1 ), .S(s4[11]) );
  ADDFX2 \intadd_41/U6  ( .A(\intadd_41/A[4] ), .B(\intadd_37/B[7] ), .CI(
        \intadd_41/n6 ), .CO(\intadd_41/n5 ), .S(\intadd_41/SUM[4] ) );
  ADDFX2 U901 ( .A(n2061), .B(\U2/Ytt[10] ), .CI(\intadd_44/n2 ), .CO(
        \intadd_44/n1 ), .S(\U2/Ytt[8] ) );
  ADDFX2 \intadd_43/U2  ( .A(n2062), .B(\U2/Xtt[10] ), .CI(\intadd_43/n2 ), 
        .CO(\intadd_43/n1 ), .S(\U2/Xtt[8] ) );
  ADDFX2 \intadd_51/U3  ( .A(\intadd_25/SUM[10] ), .B(\intadd_25/SUM[1] ), 
        .CI(\intadd_51/n3 ), .CO(\intadd_51/n2 ), .S(\U1/Xtt[1] ) );
  ADDFX2 \intadd_32/U2  ( .A(result6[11]), .B(n864), .CI(\intadd_32/n2 ), .CO(
        \intadd_32/n1 ), .S(\intadd_32/SUM[9] ) );
  ADDFX2 \intadd_30/U2  ( .A(n856), .B(n868), .CI(\intadd_30/n2 ), .CO(
        \intadd_30/n1 ), .S(s5[11]) );
  ADDFX2 \intadd_41/U5  ( .A(\intadd_41/A[5] ), .B(\intadd_37/B[8] ), .CI(
        \intadd_41/n5 ), .CO(\intadd_41/n4 ), .S(\intadd_41/SUM[5] ) );
  ADDFX2 \intadd_26/U9  ( .A(\intadd_52/n1 ), .B(\intadd_26/SUM[3] ), .CI(
        \U1/result6[13] ), .CO(\intadd_26/n8 ), .S(\U1/Ytt[3] ) );
  ADDFX2 \intadd_25/U8  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[4] ), .CI(
        \intadd_25/n8 ), .CO(\intadd_25/n7 ), .S(\U1/Xtt[4] ) );
  ADDFX2 \intadd_25/U7  ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[5] ), .CI(
        \intadd_25/n7 ), .CO(\intadd_25/n6 ), .S(\U1/Xtt[5] ) );
  OAI2BB2X1 U1666 ( .B0(n1988), .B1(n662), .A0N(n1988), .A1N(n662), .Y(n1978)
         );
  MXI2X1 U1025 ( .A(n1411), .B(n980), .S0(n1420), .Y(\U4/Yt[5] ) );
  MXI2X1 U1653 ( .A(n2579), .B(n1966), .S0(n1979), .Y(\U1/temp_xxx[2] ) );
  INVX4 U84 ( .A(n2538), .Y(n643) );
  MXI2X1 U1651 ( .A(n2346), .B(n1964), .S0(n1976), .Y(\U1/temp_xxx[3] ) );
  MXI2X1 U1365 ( .A(n732), .B(n1671), .S0(n1704), .Y(\U2/temp_x[2] ) );
  MXI2X1 U1363 ( .A(n2546), .B(n731), .S0(n1701), .Y(\U2/temp_x[3] ) );
  MXI2X1 U1361 ( .A(n1638), .B(n730), .S0(n1699), .Y(\U2/temp_x[4] ) );
  MXI2X1 U1320 ( .A(n2558), .B(n2479), .S0(n1649), .Y(\U2/temp_y[4] ) );
  AOI2BB2X1 U1317 ( .B0(n1643), .B1(n732), .A0N(n732), .A1N(n1643), .Y(n1642)
         );
  MXI2X1 U1318 ( .A(n2498), .B(n1644), .S0(n1645), .Y(\U2/temp_y[5] ) );
  MXI2X1 U1359 ( .A(n2565), .B(n745), .S0(n1697), .Y(\U2/temp_x[5] ) );
  MXI2X1 U1316 ( .A(n1641), .B(n738), .S0(n1642), .Y(\U2/temp_y[6] ) );
  MXI2X1 U1314 ( .A(n2530), .B(n739), .S0(n1639), .Y(\U2/temp_y[7] ) );
  CLKINVX3 U9 ( .A(n1221), .Y(n568) );
  AOI2BB2X1 U1567 ( .B0(n650), .B1(n1874), .A0N(n1874), .A1N(n650), .Y(n1873)
         );
  AOI2BB2X1 U1360 ( .B0(n2604), .B1(n2545), .A0N(n2545), .A1N(n2604), .Y(n1697) );
  INVX2 U28 ( .A(n1216), .Y(n587) );
  INVX2 U56 ( .A(n1198), .Y(n615) );
  CLKINVX3 U110 ( .A(n1896), .Y(n669) );
  DFFX4 \U10/temp_reg[1]  ( .D(temp4[1]), .CK(clk), .Q(temp4t[1]), .QN(n1124)
         );
  DFFHQXL \U4/U13/temp_reg[8]  ( .D(\U4/Xt[8] ), .CK(clk), .Q(result3[8]) );
  DFFHQX1 \U4/U12/temp_reg[0]  ( .D(\U4/temp7[0] ), .CK(clk), .Q(
        \U4/temp7t[0] ) );
  DFFHQX2 \U11/temp_reg[2]  ( .D(temp5[2]), .CK(clk), .Q(\U5/temp1[1] ) );
  DFFHQX1 \U1/U20/temp_reg[8]  ( .D(\U1/temp_xxx[8] ), .CK(clk), .Q(
        \U1/result5[0] ) );
  DFFHQX1 \U3/U21/temp_reg[12]  ( .D(\U3/temp10[12] ), .CK(clk), .Q(
        \U3/temp11[12] ) );
  DFFHQX1 \U1/U21/temp_reg[8]  ( .D(\U1/temp_yyy[8] ), .CK(clk), .Q(
        \U1/result6[0] ) );
  INVX4 U1800 ( .A(n2309), .Y(n2537) );
  CLKINVX3 U1801 ( .A(n2588), .Y(n769) );
  NAND2BX2 U1802 ( .AN(n775), .B(n2191), .Y(n2190) );
  INVX4 U1803 ( .A(n1931), .Y(n835) );
  NAND2X2 U1804 ( .A(n1725), .B(n2126), .Y(n2385) );
  AOI2BB2X1 U1805 ( .B0(n1279), .B1(n1273), .A0N(n1273), .A1N(n1279), .Y(n2058) );
  INVX4 U1806 ( .A(\intadd_39/n1 ), .Y(n692) );
  CLKINVX3 U1807 ( .A(n2011), .Y(n2367) );
  AOI2BB2X2 U1808 ( .B0(n1098), .B1(n1268), .A0N(n1268), .A1N(n1098), .Y(
        \intadd_39/B[7] ) );
  INVX1 U1809 ( .A(n2058), .Y(n781) );
  OAI2BB2X2 U1810 ( .B0(n1902), .B1(n1903), .A0N(n1902), .A1N(n1903), .Y(n1862) );
  INVX1 U1811 ( .A(n2002), .Y(n2379) );
  CLKINVX3 U1812 ( .A(\U5/U5/temp[5] ), .Y(n1051) );
  INVX1 U1813 ( .A(\U4/temp2[9] ), .Y(n1114) );
  INVX1 U1814 ( .A(n2795), .Y(n2703) );
  INVX1 U1815 ( .A(\U5/U5/temp[7] ), .Y(n998) );
  CLKINVX3 U1816 ( .A(\U5/U5/temp[11] ), .Y(n1021) );
  INVX1 U1817 ( .A(\intadd_37/A[6] ), .Y(n825) );
  OAI222X1 U1818 ( .A0(n636), .A1(n1140), .B0(n636), .B1(x0[1]), .C0(n1140), 
        .C1(x0[1]), .Y(n1138) );
  NAND2X1 U1819 ( .A(n1957), .B(n2346), .Y(n2466) );
  OAI222X1 U1820 ( .A0(n621), .A1(n1188), .B0(n621), .B1(x3[1]), .C0(n1188), 
        .C1(x3[1]), .Y(n1186) );
  INVX1 U1821 ( .A(\intadd_45/A[8] ), .Y(n776) );
  OAI222X1 U1822 ( .A0(n626), .A1(n1172), .B0(n626), .B1(x2[1]), .C0(n1172), 
        .C1(x2[1]), .Y(n1170) );
  OAI222X1 U1823 ( .A0(n631), .A1(n1156), .B0(n631), .B1(x1[1]), .C0(n1156), 
        .C1(x1[1]), .Y(n1154) );
  CLKINVX3 U1824 ( .A(n2380), .Y(n2536) );
  INVX1 U1825 ( .A(n1644), .Y(n2498) );
  INVX1 U1826 ( .A(n2498), .Y(n2499) );
  INVX1 U1827 ( .A(n2407), .Y(n2408) );
  INVX1 U1828 ( .A(n1715), .Y(n2400) );
  INVX1 U1829 ( .A(n1750), .Y(n2585) );
  INVX4 U1830 ( .A(n1415), .Y(n2138) );
  INVX1 U1831 ( .A(n1306), .Y(n1002) );
  CLKINVX3 U1832 ( .A(n2766), .Y(n2233) );
  CLKINVX3 U1833 ( .A(n1271), .Y(n705) );
  INVX1 U1834 ( .A(\U5/temp1[9] ), .Y(n1117) );
  MXI2X1 U1835 ( .A(n1271), .B(n705), .S0(n1246), .Y(\intadd_39/B[5] ) );
  INVX4 U1836 ( .A(n1919), .Y(n672) );
  INVX1 U1837 ( .A(n2794), .Y(n2652) );
  NOR2X1 U1838 ( .A(\U5/temp2[9] ), .B(\U5/temp1[9] ), .Y(n1294) );
  INVX1 U1839 ( .A(\U5/temp2[7] ), .Y(n1013) );
  CLKINVX3 U1840 ( .A(n738), .Y(n2133) );
  INVX1 U1841 ( .A(\U5/temp2[5] ), .Y(n1060) );
  INVX1 U1842 ( .A(\U5/temp2[6] ), .Y(n1097) );
  INVX1 U1843 ( .A(\U4/temp1[0] ), .Y(n1110) );
  INVX1 U1844 ( .A(\U5/temp2[4] ), .Y(n1096) );
  NOR2X1 U1845 ( .A(\U5/temp2[9] ), .B(n1117), .Y(n1296) );
  NAND2X1 U1846 ( .A(\U5/temp2[9] ), .B(n1117), .Y(n1297) );
  CLKINVX3 U1847 ( .A(n1244), .Y(n1098) );
  INVX1 U1848 ( .A(\intadd_47/n1 ), .Y(n804) );
  INVX1 U1849 ( .A(n2055), .Y(n780) );
  INVX1 U1850 ( .A(n2056), .Y(n779) );
  INVX1 U1851 ( .A(n1871), .Y(n652) );
  INVX1 U1852 ( .A(\U4/temp7t[2] ), .Y(n1069) );
  INVX1 U1853 ( .A(n2730), .Y(n2709) );
  INVX1 U1854 ( .A(\U5/temp5t[2] ), .Y(n1071) );
  CLKINVX3 U1855 ( .A(\U4/U6/temp[5] ), .Y(n1048) );
  INVX1 U1856 ( .A(\U4/U6/temp[7] ), .Y(n986) );
  INVX1 U1857 ( .A(n2735), .Y(n2725) );
  CLKINVX3 U1858 ( .A(\U4/U6/temp[11] ), .Y(n1020) );
  INVX1 U1859 ( .A(n2667), .Y(n2749) );
  NOR2X1 U1860 ( .A(n2667), .B(n2750), .Y(n2651) );
  CLKINVX3 U1861 ( .A(n1364), .Y(n994) );
  INVX1 U1862 ( .A(\U4/U5/temp[7] ), .Y(n974) );
  INVX1 U1863 ( .A(\U5/U6/temp[7] ), .Y(n1010) );
  NAND2X1 U1864 ( .A(n1235), .B(\U2/result2[5] ), .Y(n1252) );
  INVX1 U1865 ( .A(\U2/result2[6] ), .Y(n931) );
  NOR2X2 U1866 ( .A(n937), .B(n1253), .Y(n1235) );
  NOR2X1 U1867 ( .A(n1255), .B(n1102), .Y(n1238) );
  INVX1 U1868 ( .A(\U2/result1[8] ), .Y(n913) );
  NAND2X1 U1869 ( .A(n1236), .B(\U2/result1[5] ), .Y(n1258) );
  INVX1 U1870 ( .A(\U2/result1[6] ), .Y(n930) );
  INVX1 U1871 ( .A(\U2/result1[4] ), .Y(n936) );
  NOR2X1 U1872 ( .A(n936), .B(n1259), .Y(n1236) );
  NOR2X1 U1873 ( .A(n1261), .B(n1101), .Y(n1237) );
  XOR2X2 U1874 ( .A(n672), .B(n1920), .Y(n1922) );
  XNOR2X2 U1875 ( .A(n2589), .B(n2593), .Y(n1943) );
  CLKINVX3 U1876 ( .A(\U5/U6/temp[11] ), .Y(n1022) );
  INVX1 U1877 ( .A(\U4/U5/temp[11] ), .Y(n1019) );
  AOI2BB2X1 U1878 ( .B0(temp1t[7]), .B1(n962), .A0N(n962), .A1N(temp1t[7]), 
        .Y(n1801) );
  INVX1 U1879 ( .A(\intadd_41/B[6] ), .Y(n848) );
  OAI21X2 U1880 ( .A0(n1294), .A1(\intadd_48/n1 ), .B0(n1295), .Y(
        \intadd_38/A[6] ) );
  INVX1 U1881 ( .A(\intadd_38/A[6] ), .Y(n793) );
  INVX1 U1882 ( .A(\intadd_42/B[6] ), .Y(n803) );
  ADDFX2 U1883 ( .A(n690), .B(\intadd_33/A[5] ), .CI(\intadd_35/n3 ), .CO(
        \intadd_35/n2 ), .S(\intadd_35/SUM[8] ) );
  AOI2BB2X1 U1884 ( .B0(n738), .B1(n2131), .A0N(n727), .A1N(n738), .Y(n2517)
         );
  AOI2BB2X1 U1885 ( .B0(n2133), .B1(n2131), .A0N(n727), .A1N(n2133), .Y(n2516)
         );
  INVX1 U1886 ( .A(n1193), .Y(n608) );
  INVX1 U1887 ( .A(n1197), .Y(n614) );
  INVX1 U1888 ( .A(n1224), .Y(n572) );
  INVX1 U1889 ( .A(n1195), .Y(n611) );
  INVX1 U1890 ( .A(\intadd_37/B[2] ), .Y(n849) );
  NOR2X1 U1891 ( .A(n2568), .B(n1055), .Y(\intadd_50/CI ) );
  INVX1 U1892 ( .A(\U4/temp2[0] ), .Y(n1055) );
  OAI21XL U1893 ( .A0(n2512), .A1(n2131), .B0(n2511), .Y(n2510) );
  INVX1 U1894 ( .A(n1225), .Y(n573) );
  OAI222X1 U1895 ( .A0(n620), .A1(x3[3]), .B0(n620), .B1(n1184), .C0(x3[3]), 
        .C1(n1184), .Y(n1182) );
  MXI2X1 U1896 ( .A(n2526), .B(n2219), .S0(n1682), .Y(n1654) );
  OAI222X1 U1897 ( .A0(n635), .A1(x0[3]), .B0(n635), .B1(n1136), .C0(x0[3]), 
        .C1(n1136), .Y(n1134) );
  AOI211X1 U1898 ( .A0(n2541), .A1(n810), .B0(\intadd_47/CI ), .C0(n799), .Y(
        \intadd_38/B[0] ) );
  INVX1 U1899 ( .A(n1196), .Y(n613) );
  INVX1 U1900 ( .A(n1205), .Y(n599) );
  AOI211X2 U1901 ( .A0(n764), .A1(n1230), .B0(n2050), .C0(n719), .Y(
        \intadd_35/B[0] ) );
  INVX1 U1902 ( .A(n2552), .Y(n658) );
  OAI21X2 U1903 ( .A0(n1296), .A1(n804), .B0(n1297), .Y(\intadd_42/B[6] ) );
  OAI21X2 U1904 ( .A0(n1288), .A1(n1119), .B0(n1408), .Y(\intadd_37/A[6] ) );
  INVX1 U1905 ( .A(n1194), .Y(n610) );
  INVX1 U1906 ( .A(n1201), .Y(n592) );
  INVX1 U1907 ( .A(n1202), .Y(n594) );
  OAI222XL U1908 ( .A0(x2[4]), .A1(x5[4]), .B0(x2[4]), .B1(n597), .C0(x5[4]), 
        .C1(n597), .Y(n1203) );
  INVX1 U1909 ( .A(n1203), .Y(n596) );
  AOI222X1 U1910 ( .A0(x6[3]), .A1(x1[3]), .B0(x6[3]), .B1(n585), .C0(x1[3]), 
        .C1(n585), .Y(n1213) );
  INVX1 U1911 ( .A(n1213), .Y(n583) );
  INVX1 U1912 ( .A(n1220), .Y(n566) );
  BUFX3 U1913 ( .A(n1870), .Y(n2145) );
  OAI222X1 U1914 ( .A0(n625), .A1(x2[3]), .B0(n625), .B1(n1168), .C0(x2[3]), 
        .C1(n1168), .Y(n1166) );
  OAI222X1 U1915 ( .A0(n630), .A1(x1[3]), .B0(n630), .B1(n1152), .C0(x1[3]), 
        .C1(n1152), .Y(n1150) );
  OAI222XL U1916 ( .A0(x3[6]), .A1(x4[6]), .B0(x3[6]), .B1(n608), .C0(x4[6]), 
        .C1(n608), .Y(n1192) );
  INVX1 U1917 ( .A(n1192), .Y(n606) );
  AOI222X1 U1918 ( .A0(x1[7]), .A1(x6[7]), .B0(x1[7]), .B1(n578), .C0(x6[7]), 
        .C1(n578), .Y(n1209) );
  AOI222X1 U1919 ( .A0(x0[7]), .A1(x7[7]), .B0(x0[7]), .B1(n564), .C0(x7[7]), 
        .C1(n564), .Y(n1218) );
  INVX1 U1920 ( .A(\intadd_35/B[4] ), .Y(n699) );
  NAND2X2 U1921 ( .A(n1969), .B(n1966), .Y(n2439) );
  BUFX3 U1922 ( .A(n1698), .Y(n2604) );
  CLKINVX3 U1923 ( .A(n1641), .Y(n738) );
  INVX1 U1924 ( .A(n2558), .Y(n2479) );
  INVX1 U1925 ( .A(n1289), .Y(n1113) );
  OAI2BB1X1 U1926 ( .A0N(\intadd_28/n1 ), .A1N(n2731), .B0(n2728), .Y(n2756)
         );
  INVX1 U1927 ( .A(n2787), .Y(n2395) );
  OR2X2 U1928 ( .A(n2840), .B(n2776), .Y(n2394) );
  NOR2X1 U1929 ( .A(n1114), .B(n1118), .Y(n1288) );
  XOR2X1 U1930 ( .A(n2815), .B(n2814), .Y(n2821) );
  INVX1 U1931 ( .A(\U4/temp1[7] ), .Y(n1118) );
  INVX1 U1932 ( .A(\intadd_49/n1 ), .Y(n811) );
  CLKINVX3 U1933 ( .A(\U4/temp1[9] ), .Y(n1119) );
  INVX4 U1934 ( .A(n1412), .Y(n977) );
  CLKINVX3 U1935 ( .A(n2760), .Y(n2834) );
  NAND2X1 U1936 ( .A(n2732), .B(n2703), .Y(n2704) );
  AOI22X2 U1937 ( .A0(n999), .A1(n2457), .B0(n1302), .B1(n1002), .Y(n1300) );
  CLKINVX3 U1938 ( .A(n1302), .Y(n2137) );
  XOR2X2 U1939 ( .A(n1382), .B(n1383), .Y(n1355) );
  CLKINVX3 U1940 ( .A(n1355), .Y(n989) );
  OAI2BB1X2 U1941 ( .A0N(n2664), .A1N(n2663), .B0(n2662), .Y(n2700) );
  INVX1 U1942 ( .A(\U3/temp12[12] ), .Y(n2717) );
  NOR2X1 U1943 ( .A(n892), .B(n1251), .Y(n1231) );
  NOR2X2 U1944 ( .A(n913), .B(n1257), .Y(n1232) );
  AND2X2 U1945 ( .A(\U1/result5[0] ), .B(\U1/temp_xxxt[0] ), .Y(\intadd_25/CI ) );
  CLKINVX3 U1946 ( .A(n2015), .Y(n662) );
  INVX4 U1947 ( .A(n2014), .Y(n667) );
  BUFX12 U1948 ( .A(n1659), .Y(n2565) );
  INVX4 U1949 ( .A(n2157), .Y(n2562) );
  CLKINVX3 U1950 ( .A(n2692), .Y(n2142) );
  CLKINVX3 U1951 ( .A(n1943), .Y(n661) );
  CLKBUFX8 U1952 ( .A(n1670), .Y(n2546) );
  CLKINVX3 U1953 ( .A(n1303), .Y(n1001) );
  INVX4 U1954 ( .A(n1323), .Y(n2140) );
  INVX4 U1955 ( .A(n1327), .Y(n1008) );
  XNOR3X2 U1956 ( .A(n2144), .B(n2717), .C(n2716), .Y(n2770) );
  CLKINVX3 U1957 ( .A(n2571), .Y(n1886) );
  CLKBUFX8 U1958 ( .A(n2199), .Y(n2590) );
  INVX1 U1959 ( .A(n1989), .Y(n674) );
  INVX8 U1960 ( .A(\temp5t[0] ), .Y(n800) );
  BUFX8 U1961 ( .A(n1646), .Y(n2555) );
  CLKINVX3 U1962 ( .A(\U4/U5/temp[5] ), .Y(n1045) );
  CLKINVX3 U1963 ( .A(\U5/U6/temp[5] ), .Y(n1054) );
  INVX1 U1964 ( .A(\intadd_35/SUM[9] ), .Y(n680) );
  XOR2X1 U1965 ( .A(\intadd_33/n1 ), .B(n1516), .Y(\U3/temp9[11] ) );
  MXI2X2 U1966 ( .A(n1853), .B(n2482), .S0(n2502), .Y(\U1/temp_yyy[9] ) );
  OAI2BB1X1 U1967 ( .A0N(n1957), .A1N(n2413), .B0(n2521), .Y(n2520) );
  INVX1 U1968 ( .A(n1883), .Y(n2496) );
  INVX1 U1969 ( .A(\intadd_33/SUM[9] ), .Y(n681) );
  OAI2BB1X1 U1970 ( .A0N(n2486), .A1N(\intadd_33/n1 ), .B0(n2487), .Y(
        \U3/temp9[12] ) );
  INVX1 U1971 ( .A(n1875), .Y(n650) );
  INVX1 U1972 ( .A(\intadd_33/SUM[8] ), .Y(n682) );
  INVX1 U1973 ( .A(\intadd_33/SUM[7] ), .Y(n683) );
  INVX1 U1974 ( .A(\intadd_33/SUM[6] ), .Y(n684) );
  MXI2X1 U1975 ( .A(n1664), .B(n727), .S0(n2480), .Y(\U2/temp_x[8] ) );
  XOR2X1 U1976 ( .A(n2123), .B(n2479), .Y(n2480) );
  MXI2X2 U1977 ( .A(n1664), .B(n2131), .S0(n2485), .Y(\U2/temp_x[9] ) );
  MXI2X1 U1978 ( .A(n2530), .B(n739), .S0(n2497), .Y(\U2/temp_y[9] ) );
  MXI2X1 U1979 ( .A(n1411), .B(n980), .S0(n1413), .Y(\U4/Yt[8] ) );
  XOR2X1 U1980 ( .A(n2170), .B(n2818), .Y(\U3/Xtt[8] ) );
  XNOR2X1 U1981 ( .A(n2171), .B(n2172), .Y(\U3/Xtt[9] ) );
  OAI2BB2X2 U1982 ( .B0(n1746), .B1(n2553), .A0N(n1746), .A1N(n2553), .Y(n1659) );
  XNOR3X2 U1983 ( .A(\U3/temp9t[4] ), .B(n2606), .C(n2684), .Y(n2688) );
  CLKINVX3 U1984 ( .A(n2531), .Y(n761) );
  NAND2X1 U1985 ( .A(n1910), .B(n2550), .Y(n2180) );
  NAND2BX2 U1986 ( .AN(n1964), .B(n2345), .Y(n2344) );
  NAND2X1 U1987 ( .A(n965), .B(n1480), .Y(n2320) );
  NAND2X2 U1988 ( .A(n1725), .B(n2556), .Y(n2384) );
  NAND2X1 U1989 ( .A(n2309), .B(n1741), .Y(n2364) );
  NOR3X2 U1990 ( .A(n740), .B(n1716), .C(n1715), .Y(n1717) );
  NAND2X2 U1991 ( .A(n2130), .B(n669), .Y(n2327) );
  NAND2X2 U1992 ( .A(n1751), .B(n1750), .Y(n2403) );
  AND2X2 U1993 ( .A(n2530), .B(n730), .Y(n2484) );
  INVX1 U1994 ( .A(n763), .Y(n2201) );
  INVX1 U1995 ( .A(n2555), .Y(n734) );
  AOI2BB2X1 U1996 ( .B0(n1991), .B1(n674), .A0N(n1991), .A1N(n674), .Y(n1983)
         );
  OAI2BB2X1 U1997 ( .B0(n1996), .B1(n2587), .A0N(n1996), .A1N(n2587), .Y(n1980) );
  INVX1 U1998 ( .A(temp3t[7]), .Y(n1039) );
  INVX1 U1999 ( .A(temp2t[7]), .Y(n1037) );
  INVX1 U2000 ( .A(temp2t[6]), .Y(n1036) );
  INVX1 U2001 ( .A(temp4t[6]), .Y(n1042) );
  INVX1 U2002 ( .A(temp2t[5]), .Y(n1035) );
  INVX1 U2003 ( .A(\U4/temp5t[2] ), .Y(n1066) );
  INVX1 U2004 ( .A(\U5/temp7t[2] ), .Y(n1074) );
  CLKINVX3 U2005 ( .A(temp1t[6]), .Y(n1033) );
  INVX1 U2006 ( .A(n1893), .Y(n677) );
  MXI2X2 U2007 ( .A(n2564), .B(n760), .S0(n1827), .Y(n1679) );
  NAND2X1 U2008 ( .A(n1080), .B(temp3t[2]), .Y(n2198) );
  INVX1 U2009 ( .A(n1944), .Y(n678) );
  INVX1 U2010 ( .A(n1819), .Y(n2298) );
  NAND2X1 U2011 ( .A(temp2t[3]), .B(n1083), .Y(n2209) );
  INVX1 U2012 ( .A(n1938), .Y(n832) );
  NAND2X1 U2013 ( .A(n1903), .B(n669), .Y(n2328) );
  INVX4 U2014 ( .A(temp3t[1]), .Y(n1122) );
  XNOR2X2 U2015 ( .A(n670), .B(n1906), .Y(n1905) );
  NAND2X1 U2016 ( .A(n835), .B(n1923), .Y(n2243) );
  NAND2X1 U2017 ( .A(n1777), .B(n2358), .Y(n2265) );
  NAND2X1 U2018 ( .A(n2528), .B(n1790), .Y(n2313) );
  INVX4 U2019 ( .A(temp4t[2]), .Y(n1084) );
  NAND2X1 U2020 ( .A(n769), .B(n2548), .Y(n2254) );
  NAND2X1 U2021 ( .A(n2159), .B(n1780), .Y(n2378) );
  NAND2X1 U2022 ( .A(n1673), .B(n2561), .Y(n2175) );
  CLKINVX3 U2023 ( .A(n1909), .Y(n668) );
  INVX1 U2024 ( .A(n2159), .Y(n773) );
  NAND2X2 U2025 ( .A(n1802), .B(n962), .Y(n2160) );
  INVX1 U2026 ( .A(n1786), .Y(n770) );
  INVX1 U2027 ( .A(n1956), .Y(n837) );
  NAND2X2 U2028 ( .A(n1815), .B(n1041), .Y(n2280) );
  INVX4 U2029 ( .A(temp2t[1]), .Y(n1121) );
  INVX1 U2030 ( .A(n2128), .Y(n2574) );
  INVX4 U2031 ( .A(n1789), .Y(n754) );
  INVX4 U2032 ( .A(n2028), .Y(n673) );
  INVX1 U2033 ( .A(n775), .Y(n2192) );
  NAND2X2 U2034 ( .A(n1774), .B(n2358), .Y(n2264) );
  NAND2X2 U2035 ( .A(n1772), .B(n2588), .Y(n2353) );
  NAND2X2 U2036 ( .A(n1772), .B(n2548), .Y(n2354) );
  INVX4 U2037 ( .A(n1482), .Y(n969) );
  CLKINVX3 U2038 ( .A(n1783), .Y(n2414) );
  XOR2X2 U2039 ( .A(n1713), .B(n1721), .Y(n1719) );
  XOR2X2 U2040 ( .A(n1832), .B(n1831), .Y(n1675) );
  INVX4 U2041 ( .A(n1479), .Y(n967) );
  XOR2X2 U2042 ( .A(n772), .B(n2528), .Y(n2580) );
  INVX4 U2043 ( .A(n1777), .Y(n2293) );
  CLKBUFX8 U2044 ( .A(n2321), .Y(n1802) );
  CLKINVX3 U2045 ( .A(n2586), .Y(n767) );
  INVX8 U2046 ( .A(n2152), .Y(n2569) );
  CLKINVX3 U2047 ( .A(n2564), .Y(n760) );
  CLKINVX3 U2048 ( .A(n2539), .Y(n2240) );
  INVX4 U2049 ( .A(n1915), .Y(n2578) );
  INVX1 U2050 ( .A(temp4t[7]), .Y(n962) );
  INVX1 U2051 ( .A(n2278), .Y(n2151) );
  AOI2BB2X1 U2052 ( .B0(temp1t[9]), .B1(n1011), .A0N(n1011), .A1N(temp1t[9]), 
        .Y(n1798) );
  AOI2BB2X1 U2053 ( .B0(temp3t[9]), .B1(n1012), .A0N(n1012), .A1N(temp3t[9]), 
        .Y(n1796) );
  INVX1 U2054 ( .A(temp2t[9]), .Y(n1012) );
  INVX1 U2055 ( .A(temp4t[9]), .Y(n1011) );
  AOI22X1 U2056 ( .A0(\U5/U5/temp[4] ), .A1(n998), .B0(\U5/U5/temp[7] ), .B1(
        n1050), .Y(n2069) );
  XNOR2X1 U2057 ( .A(n1396), .B(n2069), .Y(n1379) );
  AOI22X1 U2058 ( .A0(\U5/U6/temp[6] ), .A1(n1022), .B0(\U5/U6/temp[11] ), 
        .B1(n1007), .Y(n2070) );
  XNOR2X2 U2059 ( .A(n1332), .B(n2070), .Y(n1306) );
  AOI2BB2X1 U2060 ( .B0(n1467), .B1(n963), .A0N(n963), .A1N(n1467), .Y(n2071)
         );
  MXI2X1 U2061 ( .A(n1463), .B(n968), .S0(n2071), .Y(\U4/Xt[8] ) );
  AOI2BB2X1 U2062 ( .B0(n1292), .B1(\intadd_38/n1 ), .A0N(\intadd_38/n1 ), 
        .A1N(n1292), .Y(\U5/temp5[10] ) );
  AOI2BB2X1 U2063 ( .B0(n1405), .B1(\intadd_37/n1 ), .A0N(\intadd_37/n1 ), 
        .A1N(n1405), .Y(\U4/temp5[10] ) );
  AOI22X1 U2064 ( .A0(n1306), .A1(n999), .B0(n1002), .B1(n1305), .Y(n2072) );
  MXI2X1 U2065 ( .A(n1302), .B(n2137), .S0(n2072), .Y(\U5/Yt[8] ) );
  AOI2BB2X1 U2066 ( .B0(n1272), .B1(n1273), .A0N(n1273), .A1N(n1272), .Y(
        \intadd_39/B[4] ) );
  OR2X1 U2067 ( .A(n2842), .B(n2783), .Y(n2407) );
  AOI21X1 U2068 ( .A0(n1251), .A1(n892), .B0(n1231), .Y(n2158) );
  AOI22X1 U2069 ( .A0(n980), .A1(n977), .B0(n1412), .B1(n1411), .Y(n2073) );
  XNOR2X1 U2070 ( .A(n2073), .B(n1409), .Y(\U4/Yt[9] ) );
  AOI2BB2X1 U2071 ( .B0(n973), .B1(n1469), .A0N(n1469), .A1N(n973), .Y(n2074)
         );
  MXI2X1 U2072 ( .A(n1463), .B(n968), .S0(n2074), .Y(\U4/Xt[7] ) );
  AOI2BB2X1 U2073 ( .B0(n1308), .B1(n2140), .A0N(n2140), .A1N(n1308), .Y(n2075) );
  MXI2X1 U2074 ( .A(n1302), .B(n2137), .S0(n2075), .Y(\U5/Yt[7] ) );
  AOI2BB2X1 U2075 ( .B0(n1360), .B1(n997), .A0N(n997), .A1N(n1360), .Y(n2076)
         );
  MXI2X1 U2076 ( .A(n1354), .B(n992), .S0(n2076), .Y(\U5/Xt[7] ) );
  AOI2BB2X1 U2077 ( .B0(n1266), .B1(n1267), .A0N(n1267), .A1N(n1266), .Y(
        \intadd_39/CI ) );
  AOI2BB2X1 U2078 ( .B0(n1274), .B1(n2077), .A0N(n2077), .A1N(n1274), .Y(
        \intadd_39/B[3] ) );
  INVX1 U2079 ( .A(n1248), .Y(n2077) );
  XNOR2X1 U2080 ( .A(\U3/temp10t[6] ), .B(\U3/temp10t[7] ), .Y(n2078) );
  NAND2X1 U2081 ( .A(n2078), .B(n2632), .Y(n2079) );
  OAI21XL U2082 ( .A0(n2078), .A1(n2632), .B0(n2079), .Y(n2647) );
  NAND2BX1 U2083 ( .AN(n1664), .B(n2498), .Y(n2080) );
  AOI22X4 U2084 ( .A0(n2499), .A1(n1664), .B0(n2525), .B1(n2080), .Y(n2534) );
  XNOR2X1 U2085 ( .A(n2780), .B(n2779), .Y(n2081) );
  NAND2X1 U2086 ( .A(n2081), .B(n2781), .Y(n2082) );
  OAI21XL U2087 ( .A0(n2081), .A1(n2781), .B0(n2082), .Y(n2817) );
  XNOR2X1 U2088 ( .A(\U3/temp11[1] ), .B(\U3/temp11[0] ), .Y(n2083) );
  NAND2X1 U2089 ( .A(n2083), .B(n2663), .Y(n2084) );
  OAI21X2 U2090 ( .A0(n2083), .A1(n2663), .B0(n2084), .Y(n2836) );
  NOR2BX1 U2091 ( .AN(n2839), .B(n2840), .Y(n2476) );
  AOI2BB2X1 U2092 ( .B0(n1233), .B1(\U2/result2[7] ), .A0N(\U2/result2[7] ), 
        .A1N(n1233), .Y(n2063) );
  INVX1 U2093 ( .A(n1499), .Y(n2085) );
  AOI222X4 U2094 ( .A0(n1498), .A1(n2141), .B0(n1498), .B1(n2085), .C0(n2141), 
        .C1(n2085), .Y(n1486) );
  AOI2BB2X1 U2095 ( .B0(n2163), .B1(n1435), .A0N(n1435), .A1N(n2163), .Y(n2086) );
  MXI2X1 U2096 ( .A(n985), .B(n1432), .S0(n2086), .Y(\U4/Yt[1] ) );
  AOI2BB2X1 U2097 ( .B0(n1419), .B1(n984), .A0N(n984), .A1N(n1419), .Y(n2087)
         );
  MXI2X1 U2098 ( .A(n1411), .B(n980), .S0(n2087), .Y(\U4/Yt[6] ) );
  AOI2BB2X1 U2099 ( .B0(n1362), .B1(n996), .A0N(n996), .A1N(n1362), .Y(n2088)
         );
  MXI2X1 U2100 ( .A(n1354), .B(n992), .S0(n2088), .Y(\U5/Xt[6] ) );
  INVX1 U2101 ( .A(n1463), .Y(n2089) );
  AOI21X1 U2102 ( .A0(n965), .A1(n1461), .B0(n2089), .Y(\U4/Xt[11] ) );
  INVX1 U2103 ( .A(n1302), .Y(n2090) );
  AOI21X1 U2104 ( .A0(n1001), .A1(n1300), .B0(n2090), .Y(\U5/Yt[11] ) );
  AOI2BB2X1 U2105 ( .B0(n1275), .B1(n1276), .A0N(n1276), .A1N(n1275), .Y(
        \intadd_39/B[2] ) );
  XNOR2X1 U2106 ( .A(n2779), .B(n2142), .Y(n2091) );
  NAND2X1 U2107 ( .A(n2091), .B(n2769), .Y(n2092) );
  OAI21XL U2108 ( .A0(n2091), .A1(n2769), .B0(n2092), .Y(n2778) );
  INVX1 U2109 ( .A(x4[5]), .Y(n2093) );
  AOI222X1 U2110 ( .A0(x3[5]), .A1(n1180), .B0(x3[5]), .B1(n2093), .C0(n1180), 
        .C1(n2093), .Y(n1178) );
  INVX1 U2111 ( .A(x7[5]), .Y(n2094) );
  AOI222X1 U2112 ( .A0(x0[5]), .A1(n1132), .B0(x0[5]), .B1(n2094), .C0(n1132), 
        .C1(n2094), .Y(n1130) );
  AOI22X1 U2113 ( .A0(\U4/temp2[9] ), .A1(n1118), .B0(\intadd_50/n1 ), .B1(
        n1265), .Y(n2095) );
  MXI2X1 U2114 ( .A(n1112), .B(n1263), .S0(n2095), .Y(\intadd_41/A[8] ) );
  INVX1 U2115 ( .A(x6[5]), .Y(n2096) );
  AOI222X1 U2116 ( .A0(x1[5]), .A1(n1148), .B0(x1[5]), .B1(n2096), .C0(n1148), 
        .C1(n2096), .Y(n1146) );
  INVX1 U2117 ( .A(x5[5]), .Y(n2097) );
  AOI222X1 U2118 ( .A0(x2[5]), .A1(n1164), .B0(x2[5]), .B1(n2097), .C0(n1164), 
        .C1(n2097), .Y(n1162) );
  AOI2BB2X1 U2119 ( .B0(n1191), .B1(n1175), .A0N(n1175), .A1N(n1191), .Y(
        temp4[8]) );
  AOI2BB2X1 U2120 ( .B0(n1200), .B1(n1159), .A0N(n1159), .A1N(n1200), .Y(
        temp3[8]) );
  AOI2BB2X1 U2121 ( .B0(n2552), .B1(n2522), .A0N(n2522), .A1N(n2552), .Y(n2098) );
  MXI2X1 U2122 ( .A(n654), .B(n2549), .S0(n2098), .Y(\U1/temp_yyy[6] ) );
  AOI2BB2X1 U2123 ( .B0(n1868), .B1(n1867), .A0N(n1867), .A1N(n1868), .Y(n2099) );
  MXI2X1 U2124 ( .A(n1855), .B(n2494), .S0(n2099), .Y(\U1/temp_yyy[5] ) );
  AOI2BB2X1 U2125 ( .B0(n1969), .B1(n1968), .A0N(n1968), .A1N(n1969), .Y(n2100) );
  MXI2X1 U2126 ( .A(n2579), .B(n1966), .S0(n2100), .Y(\U1/temp_xxx[6] ) );
  AOI2BB2X1 U2127 ( .B0(n1973), .B1(n2554), .A0N(n2554), .A1N(n1973), .Y(n2101) );
  MXI2X1 U2128 ( .A(n2536), .B(n2380), .S0(n2101), .Y(\U1/temp_xxx[5] ) );
  XOR2X1 U2129 ( .A(n2547), .B(n2145), .Y(n2102) );
  NAND2X1 U2130 ( .A(n2102), .B(n1871), .Y(n2103) );
  OAI21XL U2131 ( .A0(n2102), .A1(n1871), .B0(n2103), .Y(\U1/temp_yyy[4] ) );
  AOI2BB2X1 U2132 ( .B0(n639), .B1(n1975), .A0N(n1975), .A1N(n639), .Y(n2104)
         );
  MXI2X1 U2133 ( .A(n2538), .B(n643), .S0(n2104), .Y(\U1/temp_xxx[4] ) );
  AOI2BB2X1 U2134 ( .B0(n1209), .B1(n1143), .A0N(n1143), .A1N(n1209), .Y(
        temp2[8]) );
  AOI2BB2X1 U2135 ( .B0(n1218), .B1(n1127), .A0N(n1127), .A1N(n1218), .Y(
        temp1[8]) );
  AOI2BB2X1 U2136 ( .B0(n1965), .B1(n1964), .A0N(n1964), .A1N(n1965), .Y(n2105) );
  MXI2X1 U2137 ( .A(n640), .B(n1957), .S0(n2105), .Y(\U1/temp_xxx[7] ) );
  AOI2BB2X1 U2138 ( .B0(n743), .B1(n2605), .A0N(n2605), .A1N(n743), .Y(n2106)
         );
  MXI2X1 U2139 ( .A(n727), .B(n1664), .S0(n2106), .Y(\U2/temp_x[7] ) );
  XNOR2X1 U2140 ( .A(n2291), .B(n2721), .Y(n2107) );
  NAND2X1 U2141 ( .A(n2107), .B(n2722), .Y(n2108) );
  OAI21XL U2142 ( .A0(n2107), .A1(n2722), .B0(n2108), .Y(\U3/Xtt[0] ) );
  AOI2BB2X1 U2143 ( .B0(n1486), .B1(n1487), .A0N(n1487), .A1N(n1486), .Y(n2109) );
  MXI2X1 U2144 ( .A(n973), .B(n1484), .S0(n2109), .Y(\U4/Xt[1] ) );
  AOI2BB2X1 U2145 ( .B0(n1325), .B1(n1326), .A0N(n1326), .A1N(n1325), .Y(n2110) );
  MXI2X1 U2146 ( .A(n2140), .B(n1323), .S0(n2110), .Y(\U5/Yt[1] ) );
  AOI2BB2X1 U2147 ( .B0(n1377), .B1(n1378), .A0N(n1378), .A1N(n1377), .Y(n2111) );
  MXI2X1 U2148 ( .A(n997), .B(n1375), .S0(n2111), .Y(\U5/Xt[1] ) );
  AOI2BB2X1 U2149 ( .B0(n1638), .B1(n1637), .A0N(n1637), .A1N(n1638), .Y(n2112) );
  MXI2X1 U2150 ( .A(n2530), .B(n739), .S0(n2112), .Y(\U2/temp_y[8] ) );
  AOI2BB2X1 U2151 ( .B0(n985), .B1(n2470), .A0N(n2470), .A1N(n985), .Y(n2113)
         );
  MXI2X1 U2152 ( .A(n1411), .B(n980), .S0(n2113), .Y(\U4/Yt[7] ) );
  XNOR2X1 U2153 ( .A(n2809), .B(n2823), .Y(n2114) );
  NAND2X1 U2154 ( .A(n2114), .B(n2810), .Y(n2115) );
  OAI21XL U2155 ( .A0(n2114), .A1(n2810), .B0(n2115), .Y(\U3/Ytt[6] ) );
  XNOR2X1 U2156 ( .A(n2821), .B(n2839), .Y(n2116) );
  NAND2X1 U2157 ( .A(n2116), .B(n2822), .Y(n2117) );
  OAI21XL U2158 ( .A0(n2116), .A1(n2822), .B0(n2117), .Y(\U3/Xtt[6] ) );
  AOI22X1 U2159 ( .A0(n1463), .A1(n1464), .B0(n965), .B1(n968), .Y(n2118) );
  XNOR2X1 U2160 ( .A(n1461), .B(n2118), .Y(\U4/Xt[9] ) );
  XNOR2X1 U2161 ( .A(n2837), .B(n2836), .Y(n2119) );
  NAND2X1 U2162 ( .A(n2119), .B(n2838), .Y(n2120) );
  OAI21XL U2163 ( .A0(n2119), .A1(n2838), .B0(n2120), .Y(\U3/Ytt[9] ) );
  AOI22X1 U2164 ( .A0(n1001), .A1(n2137), .B0(n1303), .B1(n1302), .Y(n2121) );
  XNOR2X1 U2165 ( .A(n1300), .B(n2121), .Y(\U5/Yt[9] ) );
  AOI22X1 U2166 ( .A0(n1355), .A1(n1354), .B0(n989), .B1(n992), .Y(n2122) );
  XNOR2X1 U2167 ( .A(n1352), .B(n2122), .Y(\U5/Xt[9] ) );
  XNOR2X1 U2168 ( .A(n1254), .B(\intadd_44/n1 ), .Y(\U2/Ytt[9] ) );
  NAND2X2 U2169 ( .A(n1774), .B(n1777), .Y(n2263) );
  NAND2X2 U2170 ( .A(n1793), .B(n2548), .Y(n2253) );
  NAND2X2 U2171 ( .A(n1793), .B(n769), .Y(n2252) );
  NAND2X2 U2172 ( .A(n1357), .B(n2139), .Y(n2454) );
  OAI2BB1X4 U2173 ( .A0N(n1374), .A1N(n993), .B0(n2139), .Y(n2177) );
  INVX8 U2174 ( .A(n1476), .Y(n964) );
  INVX12 U2175 ( .A(n1484), .Y(n973) );
  INVX12 U2176 ( .A(\U4/U5/temp[1] ), .Y(n1086) );
  INVX8 U2177 ( .A(n1855), .Y(n2494) );
  AOI2BB2X1 U2178 ( .B0(n731), .B1(n1640), .A0N(n1640), .A1N(n731), .Y(n1639)
         );
  AOI2BB2X1 U2179 ( .B0(n2560), .B1(n2524), .A0N(n2524), .A1N(n2560), .Y(n1695) );
  NAND2X2 U2180 ( .A(n731), .B(n1703), .Y(n2357) );
  XOR2X4 U2181 ( .A(n1741), .B(n2331), .Y(n1739) );
  NAND2X2 U2182 ( .A(n2331), .B(n2309), .Y(n2362) );
  NAND2X2 U2183 ( .A(n2331), .B(n1741), .Y(n2363) );
  OAI2BB2X2 U2184 ( .B0(n1731), .B1(n1732), .A0N(n1731), .A1N(n1732), .Y(n1646) );
  NOR2X1 U2185 ( .A(n850), .B(n1110), .Y(\intadd_46/CI ) );
  NAND2X4 U2186 ( .A(n1738), .B(n2531), .Y(n2299) );
  MXI2X1 U2187 ( .A(n1853), .B(n2482), .S0(n1860), .Y(\U1/temp_yyy[7] ) );
  MX2X1 U2188 ( .A(n2482), .B(n1853), .S0(n2458), .Y(\U1/temp_yyy[8] ) );
  XOR2X2 U2189 ( .A(n2533), .B(n2547), .Y(n2458) );
  XNOR2X2 U2190 ( .A(n1937), .B(n1939), .Y(n1885) );
  BUFX16 U2191 ( .A(n1733), .Y(n2147) );
  NAND2X4 U2192 ( .A(n1706), .B(n1705), .Y(n2337) );
  NAND2X4 U2193 ( .A(n1676), .B(n1673), .Y(n2174) );
  INVX16 U2194 ( .A(n2127), .Y(n664) );
  INVX16 U2195 ( .A(n1964), .Y(n2346) );
  NAND2X4 U2196 ( .A(n2380), .B(n646), .Y(n2431) );
  BUFX16 U2197 ( .A(n1833), .Y(n2539) );
  BUFX16 U2198 ( .A(n1849), .Y(n2542) );
  BUFX16 U2199 ( .A(n2258), .Y(n1706) );
  NAND2X2 U2200 ( .A(n2210), .B(n2688), .Y(n2221) );
  OAI2BB1X4 U2201 ( .A0N(n2383), .A1N(n2721), .B0(n2291), .Y(n2381) );
  NAND2X2 U2202 ( .A(\U3/temp11[0] ), .B(\U3/temp9t[0] ), .Y(n2669) );
  NAND2X4 U2203 ( .A(n1715), .B(n1750), .Y(n2404) );
  AOI2BB2X4 U2204 ( .B0(n2606), .B1(n2717), .A0N(n2716), .A1N(n2715), .Y(n2842) );
  INVX4 U2205 ( .A(n2813), .Y(n2719) );
  XNOR3X2 U2206 ( .A(\U3/temp12[0] ), .B(n2606), .C(n2680), .Y(n2813) );
  AND3X4 U2207 ( .A(n2450), .B(n2452), .C(n2451), .Y(n2123) );
  OAI2BB2X4 U2208 ( .B0(n1891), .B1(n671), .A0N(n1891), .A1N(n671), .Y(n1867)
         );
  XNOR2X4 U2209 ( .A(n1844), .B(n1841), .Y(n2124) );
  XOR2X4 U2210 ( .A(n2038), .B(n2573), .Y(n2125) );
  XNOR2X4 U2211 ( .A(n1716), .B(n1762), .Y(n1664) );
  XNOR2X4 U2212 ( .A(n1766), .B(n1767), .Y(n2126) );
  XOR2X4 U2213 ( .A(n1774), .B(n1775), .Y(n1732) );
  XOR2X4 U2214 ( .A(n2021), .B(n1918), .Y(n2127) );
  XOR2X4 U2215 ( .A(n1795), .B(n1788), .Y(n2434) );
  AOI2BB2X4 U2216 ( .B0(n1726), .B1(n2562), .A0N(n1726), .A1N(n2562), .Y(n1671) );
  XOR2X2 U2217 ( .A(n1945), .B(n1946), .Y(n1893) );
  OAI2BB2X4 U2218 ( .B0(n1722), .B1(n2563), .A0N(n1722), .A1N(n2563), .Y(n1638) );
  XNOR2X4 U2219 ( .A(n2029), .B(n1806), .Y(n1928) );
  INVX1 U2220 ( .A(n2689), .Y(n2720) );
  XOR2X1 U2221 ( .A(n2129), .B(n2401), .Y(n2497) );
  CLKINVX3 U2222 ( .A(n1358), .Y(n2139) );
  BUFX12 U2223 ( .A(n1804), .Y(n2128) );
  XOR2X2 U2224 ( .A(n1840), .B(n1820), .Y(n1804) );
  MX2X4 U2225 ( .A(n2519), .B(n2518), .S0(n2534), .Y(\U2/temp_x[10] ) );
  BUFX16 U2226 ( .A(n1635), .Y(n2129) );
  BUFX16 U2227 ( .A(n1908), .Y(n2130) );
  BUFX12 U2228 ( .A(n1633), .Y(n2530) );
  INVX8 U2229 ( .A(n1664), .Y(n2131) );
  BUFX12 U2230 ( .A(n2374), .Y(n1853) );
  INVX12 U2231 ( .A(n1957), .Y(n640) );
  XOR2X1 U2232 ( .A(n2827), .B(n2805), .Y(\U3/Ytt[8] ) );
  INVX4 U2233 ( .A(n2722), .Y(n2383) );
  ADDFX2 U2234 ( .A(\intadd_33/A[1] ), .B(\intadd_35/B[4] ), .CI(
        \intadd_35/n7 ), .CO(\intadd_35/n6 ), .S(\intadd_35/SUM[4] ) );
  ADDFX2 U2235 ( .A(\intadd_33/A[0] ), .B(\intadd_35/B[3] ), .CI(
        \intadd_35/n8 ), .CO(\intadd_35/n7 ), .S(\intadd_35/SUM[3] ) );
  ADDFX2 U2236 ( .A(\U1/result5[13] ), .B(\intadd_25/SUM[2] ), .CI(
        \intadd_51/n2 ), .CO(\intadd_51/n1 ), .S(\U1/Xtt[2] ) );
  OAI2BB1X2 U2237 ( .A0N(n2628), .A1N(n2630), .B0(n2627), .Y(n2663) );
  INVX4 U2238 ( .A(n2647), .Y(n2750) );
  ADDFX2 U2239 ( .A(\U1/result5[0] ), .B(\U1/result5[13] ), .CI(
        \intadd_25/n14 ), .CO(\intadd_25/n13 ), .S(\intadd_25/SUM[7] ) );
  INVX2 U2240 ( .A(n1222), .Y(n569) );
  INVX2 U2241 ( .A(n1204), .Y(n597) );
  INVX20 U2242 ( .A(n2606), .Y(n2144) );
  INVX4 U2243 ( .A(temp2t[3]), .Y(n1081) );
  INVX8 U2244 ( .A(\U3/temp11[12] ), .Y(n2606) );
  INVX2 U2245 ( .A(n1207), .Y(n601) );
  NAND2BX2 U2246 ( .AN(n2482), .B(n2134), .Y(n2447) );
  NAND2BX1 U2247 ( .AN(n2482), .B(n2494), .Y(n2493) );
  NAND2BX1 U2248 ( .AN(n1853), .B(n2547), .Y(n2481) );
  INVX4 U2249 ( .A(n2401), .Y(n2545) );
  NAND2BX1 U2250 ( .AN(n2536), .B(n640), .Y(n2515) );
  NAND2X1 U2251 ( .A(n640), .B(n643), .Y(n2492) );
  XOR2X1 U2252 ( .A(n2808), .B(n2807), .Y(\U3/Ytt[7] ) );
  AND2X2 U2253 ( .A(n2787), .B(n2778), .Y(n2396) );
  INVX1 U2254 ( .A(n2841), .Y(n2478) );
  CLKBUFX8 U2255 ( .A(n2375), .Y(n2840) );
  ADDFX2 U2256 ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[10] ), .CI(
        \intadd_26/n2 ), .CO(\U1/Ytt[11] ), .S(\U1/Ytt[10] ) );
  ADDFX2 U2257 ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[9] ), .CI(
        \intadd_26/n3 ), .CO(\intadd_26/n2 ), .S(\U1/Ytt[9] ) );
  NOR2X1 U2258 ( .A(n2232), .B(n2842), .Y(n2419) );
  INVX4 U2259 ( .A(n2829), .Y(n2830) );
  INVX1 U2260 ( .A(n2811), .Y(n2815) );
  INVX1 U2261 ( .A(n2817), .Y(n2416) );
  INVX4 U2262 ( .A(n1747), .Y(n2132) );
  INVX1 U2263 ( .A(n2806), .Y(n2804) );
  INVX1 U2264 ( .A(n2809), .Y(n2800) );
  NAND2X1 U2265 ( .A(n2136), .B(n2842), .Y(n2768) );
  ADDFX2 U2266 ( .A(\intadd_51/n1 ), .B(\intadd_25/SUM[3] ), .CI(
        \U1/result5[13] ), .CO(\intadd_25/n8 ), .S(\U1/Xtt[3] ) );
  INVX1 U2267 ( .A(n2796), .Y(n2799) );
  OAI21XL U2268 ( .A0(x5[8]), .A1(x2[8]), .B0(n1200), .Y(n1199) );
  OAI21X2 U2269 ( .A0(n1115), .A1(n1097), .B0(n705), .Y(n1519) );
  INVX1 U2270 ( .A(n2755), .Y(n2744) );
  ADDFX2 U2271 ( .A(\intadd_26/SUM[10] ), .B(\intadd_26/SUM[1] ), .CI(
        \intadd_52/n3 ), .CO(\intadd_52/n2 ), .S(\U1/Ytt[1] ) );
  CLKINVX3 U2272 ( .A(n1219), .Y(n564) );
  AOI2BB2X2 U2273 ( .B0(n2144), .B1(\U3/temp12[0] ), .A0N(n2680), .A1N(n2678), 
        .Y(n2696) );
  ADDFX2 U2274 ( .A(\U1/result6[2] ), .B(\U1/result6[13] ), .CI(
        \intadd_26/n12 ), .CO(\intadd_26/SUM[10] ), .S(\intadd_26/SUM[9] ) );
  AOI2BB2X2 U2275 ( .B0(n2144), .B1(\U3/temp9t[8] ), .A0N(n2681), .A1N(n2676), 
        .Y(n2679) );
  INVX4 U2276 ( .A(n1277), .Y(n720) );
  AND2X2 U2277 ( .A(\U3/temp12[12] ), .B(n2144), .Y(n2715) );
  CLKINVX3 U2278 ( .A(n1206), .Y(n600) );
  INVX4 U2279 ( .A(temp2t[2]), .Y(n1080) );
  INVX4 U2280 ( .A(n1959), .Y(n2592) );
  MXI2X2 U2281 ( .A(n640), .B(n1957), .S0(n2488), .Y(\U1/temp_xxx[8] ) );
  BUFX3 U2282 ( .A(n2523), .Y(n2605) );
  INVX16 U2283 ( .A(n2530), .Y(n739) );
  INVX20 U2284 ( .A(n2308), .Y(n2522) );
  XOR2X2 U2285 ( .A(n2477), .B(n2478), .Y(n2843) );
  MXI2X1 U2286 ( .A(n1651), .B(n743), .S0(n1652), .Y(\U2/temp_y[3] ) );
  AOI2BB2X1 U2287 ( .B0(n1653), .B1(n1654), .A0N(n1654), .A1N(n1653), .Y(n1652) );
  INVX4 U2288 ( .A(n1638), .Y(n730) );
  BUFX12 U2289 ( .A(n1648), .Y(n2558) );
  XOR2X1 U2290 ( .A(n2816), .B(n2782), .Y(\U3/Xtt[5] ) );
  XOR2X2 U2291 ( .A(n2333), .B(n2013), .Y(n2012) );
  INVX16 U2292 ( .A(n1651), .Y(n743) );
  XOR2X1 U2293 ( .A(n2785), .B(n2784), .Y(\U3/Xtt[4] ) );
  INVX4 U2294 ( .A(n2838), .Y(n2831) );
  XOR2X1 U2295 ( .A(n2789), .B(n2788), .Y(\U3/Xtt[3] ) );
  INVX20 U2296 ( .A(n1655), .Y(n744) );
  XOR2X1 U2297 ( .A(n2792), .B(n2791), .Y(\U3/Xtt[2] ) );
  INVX8 U2298 ( .A(n2436), .Y(n1655) );
  XOR2X1 U2299 ( .A(n2723), .B(n2777), .Y(\U3/Xtt[1] ) );
  INVX16 U2300 ( .A(n2544), .Y(n2134) );
  XOR2X1 U2301 ( .A(n2840), .B(n2776), .Y(n2723) );
  INVX4 U2302 ( .A(n2000), .Y(n2325) );
  XOR2X1 U2303 ( .A(n2798), .B(n2751), .Y(\U3/Ytt[5] ) );
  XOR2X1 U2304 ( .A(n2754), .B(n2753), .Y(\U3/Ytt[4] ) );
  INVX4 U2305 ( .A(n2579), .Y(n1966) );
  NAND2X1 U2306 ( .A(n2291), .B(n2839), .Y(n2426) );
  NAND2BX1 U2307 ( .AN(n2291), .B(n2842), .Y(n2425) );
  XNOR3X2 U2308 ( .A(n2839), .B(n2233), .C(n2295), .Y(n2375) );
  BUFX12 U2309 ( .A(n1972), .Y(n2554) );
  XOR2X1 U2310 ( .A(n2758), .B(n2757), .Y(\U3/Ytt[3] ) );
  BUFX20 U2311 ( .A(n1728), .Y(n2553) );
  BUFX12 U2312 ( .A(n2368), .Y(n1748) );
  BUFX12 U2313 ( .A(n1745), .Y(n2156) );
  INVX4 U2314 ( .A(n2580), .Y(n2135) );
  AND2X2 U2315 ( .A(n2756), .B(n2755), .Y(n2743) );
  NAND2BX1 U2316 ( .AN(n2821), .B(n2839), .Y(n2418) );
  NAND2X1 U2317 ( .A(n2821), .B(n2842), .Y(n2417) );
  NAND2X1 U2318 ( .A(n2825), .B(\intadd_28/n1 ), .Y(n2826) );
  ADDFX2 U2319 ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[5] ), .CI(
        \intadd_26/n7 ), .CO(\intadd_26/n6 ), .S(\U1/Ytt[5] ) );
  NAND2X1 U2320 ( .A(n2800), .B(\intadd_28/n1 ), .Y(n2801) );
  BUFX12 U2321 ( .A(n1737), .Y(n2531) );
  NOR2X2 U2322 ( .A(n2842), .B(n2233), .Y(n2246) );
  ADDFX2 U2323 ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[4] ), .CI(
        \intadd_26/n8 ), .CO(\intadd_26/n7 ), .S(\U1/Ytt[4] ) );
  OAI21X2 U2324 ( .A0(\U5/temp2[6] ), .A1(\U5/temp1[6] ), .B0(n1519), .Y(n1269) );
  ADDFX2 U2325 ( .A(\U1/result6[13] ), .B(\intadd_26/SUM[2] ), .CI(
        \intadd_52/n2 ), .CO(\intadd_52/n1 ), .S(\U1/Ytt[2] ) );
  INVX8 U2326 ( .A(n2770), .Y(n2136) );
  NAND2X2 U2327 ( .A(n2719), .B(n2812), .Y(n2227) );
  BUFX20 U2328 ( .A(n1679), .Y(n2566) );
  BUFX12 U2329 ( .A(n1675), .Y(n2561) );
  AOI22X4 U2330 ( .A0(n1832), .A1(n2239), .B0(n1838), .B1(n2539), .Y(n1834) );
  INVX8 U2331 ( .A(n2290), .Y(n2588) );
  AND2X2 U2332 ( .A(\intadd_26/SUM[8] ), .B(n2303), .Y(\intadd_52/B[0] ) );
  INVX8 U2333 ( .A(n1803), .Y(n768) );
  XOR2X1 U2334 ( .A(n1231), .B(\U2/result2[9] ), .Y(n2061) );
  INVX4 U2335 ( .A(n1927), .Y(n833) );
  INVX8 U2336 ( .A(n1488), .Y(n2141) );
  OAI222X4 U2337 ( .A0(x0[4]), .A1(x7[4]), .B0(x0[4]), .B1(n569), .C0(x7[4]), 
        .C1(n569), .Y(n1221) );
  NAND2X2 U2338 ( .A(n1234), .B(\U2/result1[7] ), .Y(n1257) );
  NAND2X2 U2339 ( .A(n1233), .B(\U2/result2[7] ), .Y(n1251) );
  XOR2X4 U2340 ( .A(n2039), .B(n1840), .Y(n1940) );
  XOR2X4 U2341 ( .A(n2041), .B(n1844), .Y(n1956) );
  INVX4 U2342 ( .A(n1230), .Y(n801) );
  BUFX12 U2343 ( .A(n1282), .Y(n2551) );
  INVX8 U2344 ( .A(\temp7t[0] ), .Y(n850) );
  CLKINVX8 U2345 ( .A(n2541), .Y(n851) );
  CLKINVX3 U2346 ( .A(n1821), .Y(n2143) );
  BUFX12 U2347 ( .A(\temp6t[0] ), .Y(n2568) );
  BUFX20 U2348 ( .A(\temp8t[0] ), .Y(n2541) );
  AOI2BB2X4 U2349 ( .B0(temp2t[4]), .B1(temp3t[4]), .A0N(temp3t[4]), .A1N(
        temp2t[4]), .Y(n1840) );
  INVX1 U2350 ( .A(\U5/temp2[2] ), .Y(n1125) );
  INVX1 U2351 ( .A(\intadd_35/SUM[7] ), .Y(n686) );
  AND2X2 U2352 ( .A(n1802), .B(temp1t[7]), .Y(n2372) );
  INVX1 U2353 ( .A(\intadd_35/SUM[6] ), .Y(n687) );
  INVX1 U2354 ( .A(\intadd_35/SUM[8] ), .Y(n685) );
  AOI2BB2X1 U2355 ( .B0(\U5/temp1[1] ), .B1(\U5/temp2[1] ), .A0N(\U5/temp2[1] ), .A1N(\U5/temp1[1] ), .Y(n1267) );
  INVX1 U2356 ( .A(\U5/temp2[1] ), .Y(n1099) );
  NAND2X1 U2357 ( .A(n1034), .B(temp3t[4]), .Y(n2257) );
  NAND2BX1 U2358 ( .AN(\U3/temp12[12] ), .B(\U3/temp10t[2] ), .Y(n2611) );
  NAND2BX1 U2359 ( .AN(\U3/temp10t[2] ), .B(\U3/temp12[12] ), .Y(n2612) );
  XNOR3X2 U2360 ( .A(\U3/temp10t[3] ), .B(n2638), .C(n2637), .Y(n2708) );
  NAND2BX1 U2361 ( .AN(\U3/temp10t[3] ), .B(\U3/temp10t[4] ), .Y(n2615) );
  NAND2BX1 U2362 ( .AN(\U3/temp10t[3] ), .B(\U3/temp10t[2] ), .Y(n2614) );
  NAND2BX1 U2363 ( .AN(\U3/temp10t[2] ), .B(\U3/temp10t[3] ), .Y(n2613) );
  AOI2BB2X1 U2364 ( .B0(temp1t[5]), .B1(n1041), .A0N(n1041), .A1N(temp1t[5]), 
        .Y(n1821) );
  NAND2X2 U2365 ( .A(n1815), .B(temp1t[5]), .Y(n2279) );
  INVX1 U2366 ( .A(\U5/U5/temp[6] ), .Y(n995) );
  INVX1 U2367 ( .A(\U5/U6/temp[6] ), .Y(n1007) );
  INVX1 U2368 ( .A(\U4/U5/temp[6] ), .Y(n971) );
  INVX4 U2369 ( .A(n1421), .Y(n982) );
  AOI2BB2X2 U2370 ( .B0(\intadd_45/n1 ), .B1(n1284), .A0N(n1284), .A1N(
        \intadd_45/n1 ), .Y(n2052) );
  INVX4 U2371 ( .A(\intadd_45/n1 ), .Y(n694) );
  AOI22X4 U2372 ( .A0(n2560), .A1(n726), .B0(n1668), .B1(n728), .Y(n1666) );
  NAND2BX4 U2373 ( .AN(n1838), .B(n2240), .Y(n2239) );
  BUFX12 U2374 ( .A(n1677), .Y(n2146) );
  XOR2X2 U2375 ( .A(n1830), .B(n1831), .Y(n1677) );
  XNOR3X2 U2376 ( .A(\U3/temp11[0] ), .B(\U3/temp10t[9] ), .C(n2630), .Y(n2795) );
  XOR2X4 U2377 ( .A(n1995), .B(n662), .Y(n1994) );
  INVX12 U2378 ( .A(temp1t[2]), .Y(n1079) );
  MXI2X1 U2379 ( .A(n1655), .B(n744), .S0(n1695), .Y(\U2/temp_x[6] ) );
  XOR2X4 U2380 ( .A(n1896), .B(n2130), .Y(n1907) );
  OAI2BB1X4 U2381 ( .A0N(n1411), .A1N(n2470), .B0(n985), .Y(n2489) );
  XNOR2X4 U2382 ( .A(n1444), .B(n2282), .Y(n1432) );
  NAND2X4 U2383 ( .A(n2539), .B(n2576), .Y(n2154) );
  INVX8 U2384 ( .A(n1997), .Y(n676) );
  NOR2X4 U2385 ( .A(n1997), .B(n2587), .Y(n2596) );
  NAND2BX1 U2386 ( .AN(\U3/temp12[1] ), .B(\U3/temp10t[1] ), .Y(n2610) );
  NAND2X1 U2387 ( .A(\U3/temp12[1] ), .B(n2608), .Y(n2609) );
  AOI2BB2X4 U2388 ( .B0(n775), .B1(n1829), .A0N(n775), .A1N(n1829), .Y(n1827)
         );
  INVX8 U2389 ( .A(n1672), .Y(n725) );
  MXI2X1 U2390 ( .A(n2544), .B(n2134), .S0(n1873), .Y(\U1/temp_yyy[3] ) );
  AOI2BB2X1 U2391 ( .B0(n2134), .B1(n2535), .A0N(n2134), .A1N(n2535), .Y(n1860) );
  NAND2X1 U2392 ( .A(temp2t[5]), .B(n1038), .Y(n2148) );
  NAND2X2 U2393 ( .A(temp2t[5]), .B(n1816), .Y(n2149) );
  NAND2X2 U2394 ( .A(n1038), .B(n1816), .Y(n2150) );
  AND3X4 U2395 ( .A(n2148), .B(n2149), .C(n2150), .Y(n1809) );
  XOR2X2 U2396 ( .A(n1809), .B(n2342), .Y(n2341) );
  XOR2X4 U2397 ( .A(n2276), .B(n1799), .Y(n2370) );
  NAND2BX4 U2398 ( .AN(n2570), .B(n1955), .Y(n2152) );
  INVX12 U2399 ( .A(n1688), .Y(n752) );
  AOI22X4 U2400 ( .A0(n1809), .A1(n2277), .B0(n2151), .B1(n1036), .Y(n2276) );
  XNOR2X4 U2401 ( .A(n1907), .B(n1903), .Y(n1855) );
  BUFX16 U2402 ( .A(n1828), .Y(n2564) );
  OR2X2 U2403 ( .A(n2157), .B(n2553), .Y(n2332) );
  XNOR2X4 U2404 ( .A(n1816), .B(n2298), .Y(n2297) );
  XOR2X4 U2405 ( .A(n1843), .B(n1846), .Y(n2206) );
  MXI2X1 U2406 ( .A(\intadd_35/n1 ), .B(n679), .S0(n1516), .Y(\U3/temp10[11] )
         );
  ADDFX2 U2407 ( .A(n691), .B(n2052), .CI(\intadd_33/n2 ), .CO(\intadd_33/n1 ), 
        .S(\intadd_33/SUM[9] ) );
  INVX4 U2408 ( .A(n2052), .Y(n688) );
  XOR2X4 U2409 ( .A(n1750), .B(n1757), .Y(n1756) );
  XOR2X4 U2410 ( .A(n2582), .B(n1806), .Y(n2358) );
  INVX8 U2411 ( .A(n1687), .Y(n748) );
  NAND2X4 U2412 ( .A(n637), .B(n2579), .Y(n2188) );
  ADDFX2 U2413 ( .A(\intadd_26/SUM[9] ), .B(\intadd_52/B[0] ), .CI(
        \intadd_26/SUM[0] ), .CO(\intadd_52/n3 ), .S(\U1/Ytt[0] ) );
  OAI2BB1X4 U2414 ( .A0N(n1953), .A1N(n2569), .B0(n1954), .Y(n2042) );
  INVX20 U2415 ( .A(n2570), .Y(n1240) );
  XOR2X1 U2416 ( .A(n2820), .B(n2819), .Y(\U3/Xtt[7] ) );
  XOR2X4 U2417 ( .A(n1915), .B(n1916), .Y(n1899) );
  AOI21X4 U2418 ( .A0(n2549), .A1(n1882), .B0(n1853), .Y(\U1/temp_yyy[11] ) );
  NAND2X4 U2419 ( .A(n1738), .B(n758), .Y(n2300) );
  OAI21X1 U2420 ( .A0(\U5/temp2[0] ), .A1(n787), .B0(n1518), .Y(n1281) );
  OAI22X2 U2421 ( .A0(n678), .A1(n2584), .B0(n1826), .B1(n1944), .Y(n1992) );
  NAND2X4 U2422 ( .A(n2539), .B(n1830), .Y(n2153) );
  NAND2X4 U2423 ( .A(n1830), .B(n2576), .Y(n2155) );
  AND3X4 U2424 ( .A(n2153), .B(n2154), .C(n2155), .Y(n1824) );
  INVX8 U2425 ( .A(n2124), .Y(n2212) );
  XOR2X1 U2426 ( .A(n2765), .B(n2764), .Y(n2783) );
  XOR2X4 U2427 ( .A(n1882), .B(n2496), .Y(\U1/temp_yyy[10] ) );
  NAND2X4 U2428 ( .A(n2552), .B(n1878), .Y(n2182) );
  XOR2X4 U2429 ( .A(n1951), .B(n1952), .Y(n1946) );
  NAND2X4 U2430 ( .A(n2568), .B(\temp7t[0] ), .Y(n2043) );
  XOR2X4 U2431 ( .A(n1938), .B(n1936), .Y(n1939) );
  XOR2X4 U2432 ( .A(n1776), .B(n1775), .Y(n1728) );
  ADDFHX4 U2433 ( .A(n691), .B(n695), .CI(\intadd_33/n3 ), .CO(\intadd_33/n2 ), 
        .S(\intadd_33/SUM[8] ) );
  NOR2X2 U2434 ( .A(\intadd_35/A[2] ), .B(n765), .Y(n1228) );
  AOI22X2 U2435 ( .A0(n2567), .A1(n801), .B0(n1230), .B1(n724), .Y(
        \intadd_45/B[0] ) );
  AOI22X2 U2436 ( .A0(\U5/temp2[0] ), .A1(n810), .B0(\U5/temp1[0] ), .B1(n852), 
        .Y(n1230) );
  OR2X4 U2437 ( .A(n1744), .B(n2219), .Y(n2369) );
  XOR2X4 U2438 ( .A(n2572), .B(n1948), .Y(n2571) );
  XOR2X4 U2439 ( .A(n1956), .B(n1950), .Y(n1948) );
  XNOR2X4 U2440 ( .A(n2556), .B(n1755), .Y(n1754) );
  NAND2X4 U2441 ( .A(n1698), .B(n2401), .Y(n2420) );
  XOR2X4 U2442 ( .A(n2553), .B(n733), .Y(n1726) );
  NAND2X2 U2443 ( .A(n732), .B(n1705), .Y(n2339) );
  XOR2X4 U2444 ( .A(n762), .B(n2147), .Y(n1731) );
  NAND2X2 U2445 ( .A(n1706), .B(n732), .Y(n2338) );
  XOR2X4 U2446 ( .A(n1927), .B(n1928), .Y(n1935) );
  XOR2X4 U2447 ( .A(n1793), .B(n1773), .Y(n1747) );
  NAND2X4 U2448 ( .A(n1655), .B(n737), .Y(n2440) );
  BUFX16 U2449 ( .A(n1661), .Y(n2529) );
  XOR2X4 U2450 ( .A(n1752), .B(n2435), .Y(n2436) );
  XNOR2X4 U2451 ( .A(n1732), .B(n1753), .Y(n1752) );
  CLKINVX3 U2452 ( .A(n850), .Y(n2602) );
  NAND2X4 U2453 ( .A(n1870), .B(n652), .Y(n2260) );
  NAND2X4 U2454 ( .A(n1870), .B(n2547), .Y(n2261) );
  NAND2X4 U2455 ( .A(n1878), .B(n1877), .Y(n2183) );
  XOR2X4 U2456 ( .A(n1940), .B(n2125), .Y(n1949) );
  NAND2X4 U2457 ( .A(n1655), .B(n1658), .Y(n2441) );
  AOI21X4 U2458 ( .A0(n2413), .A1(n2514), .B0(n640), .Y(\U1/temp_xxx[11] ) );
  MXI2X4 U2459 ( .A(n2530), .B(n739), .S0(n1666), .Y(\U2/temp_y[10] ) );
  AOI2BB2X1 U2460 ( .B0(n2555), .B1(n1647), .A0N(n1647), .A1N(n2555), .Y(n1645) );
  XOR2X4 U2461 ( .A(n1748), .B(n2132), .Y(n1746) );
  OAI2BB1X4 U2462 ( .A0N(n2565), .A1N(n746), .B0(n2317), .Y(n2316) );
  NAND2X4 U2463 ( .A(n2531), .B(n758), .Y(n2301) );
  XOR2X4 U2464 ( .A(n768), .B(n2128), .Y(n1837) );
  ADDFHX4 U2465 ( .A(n690), .B(\intadd_33/A[6] ), .CI(\intadd_35/n2 ), .CO(
        \intadd_35/n1 ), .S(\intadd_35/SUM[9] ) );
  INVX4 U2466 ( .A(\intadd_45/SUM[2] ), .Y(n719) );
  OAI2BB2X4 U2467 ( .B0(n1743), .B1(n2526), .A0N(n1743), .A1N(n2526), .Y(n1686) );
  XOR2X4 U2468 ( .A(n1744), .B(n2156), .Y(n1743) );
  XOR2X4 U2469 ( .A(n766), .B(n2539), .Y(n1831) );
  OR2X4 U2470 ( .A(n748), .B(n1730), .Y(n2228) );
  OAI2BB1X4 U2471 ( .A0N(n2694), .A1N(n2688), .B0(n2687), .Y(n2214) );
  OAI222X4 U2472 ( .A0(x2[6]), .A1(x5[6]), .B0(x2[6]), .B1(n594), .C0(x5[6]), 
        .C1(n594), .Y(n1201) );
  AOI222X4 U2473 ( .A0(x5[5]), .A1(x2[5]), .B0(x5[5]), .B1(n596), .C0(x2[5]), 
        .C1(n596), .Y(n1202) );
  AOI222X4 U2474 ( .A0(x2[1]), .A1(x5[1]), .B0(x2[1]), .B1(n601), .C0(x5[1]), 
        .C1(n601), .Y(n1206) );
  AOI222X4 U2475 ( .A0(x2[7]), .A1(x5[7]), .B0(x2[7]), .B1(n592), .C0(x5[7]), 
        .C1(n592), .Y(n1200) );
  AOI222X4 U2476 ( .A0(x7[5]), .A1(x0[5]), .B0(x7[5]), .B1(n568), .C0(x0[5]), 
        .C1(n568), .Y(n1220) );
  AOI222X4 U2477 ( .A0(x0[1]), .A1(x7[1]), .B0(x0[1]), .B1(n573), .C0(x7[1]), 
        .C1(n573), .Y(n1224) );
  AOI222X4 U2478 ( .A0(x7[3]), .A1(x0[3]), .B0(x7[3]), .B1(n571), .C0(x0[3]), 
        .C1(n571), .Y(n1222) );
  OAI222X4 U2479 ( .A0(n570), .A1(x7[2]), .B0(n570), .B1(n1138), .C0(x7[2]), 
        .C1(n1138), .Y(n1136) );
  OAI222X4 U2480 ( .A0(n598), .A1(x5[2]), .B0(n598), .B1(n1170), .C0(x5[2]), 
        .C1(n1170), .Y(n1168) );
  OAI222X4 U2481 ( .A0(n609), .A1(x4[4]), .B0(n609), .B1(n1182), .C0(x4[4]), 
        .C1(n1182), .Y(n1180) );
  OAI222X4 U2482 ( .A0(n581), .A1(x6[4]), .B0(n581), .B1(n1150), .C0(x6[4]), 
        .C1(n1150), .Y(n1148) );
  OAI222X4 U2483 ( .A0(x3[4]), .A1(x4[4]), .B0(x3[4]), .B1(n611), .C0(x4[4]), 
        .C1(n611), .Y(n1194) );
  NAND2X2 U2484 ( .A(n2834), .B(n2740), .Y(n2741) );
  AND2X4 U2485 ( .A(n2806), .B(n2659), .Y(n2710) );
  AOI2BB2X2 U2486 ( .B0(n2709), .B1(n2657), .A0N(n2707), .A1N(n2643), .Y(n2733) );
  OAI222X4 U2487 ( .A0(x1[6]), .A1(x6[6]), .B0(x1[6]), .B1(n580), .C0(x6[6]), 
        .C1(n580), .Y(n1210) );
  OAI222X4 U2488 ( .A0(x1[2]), .A1(x6[2]), .B0(x1[2]), .B1(n586), .C0(x6[2]), 
        .C1(n586), .Y(n1214) );
  XNOR2X4 U2489 ( .A(n1335), .B(n1336), .Y(n1323) );
  NOR2BX2 U2490 ( .AN(\intadd_45/B[0] ), .B(n764), .Y(n2050) );
  NOR2X2 U2491 ( .A(n2383), .B(n2721), .Y(n2382) );
  NAND2X2 U2492 ( .A(n2840), .B(n2776), .Y(n2393) );
  NAND2X2 U2493 ( .A(n2213), .B(n2689), .Y(n2220) );
  NAND2BX4 U2494 ( .AN(\U4/temp5t[0] ), .B(\U4/U5/temp[0] ), .Y(n1507) );
  NAND2X2 U2495 ( .A(n654), .B(n658), .Y(n2348) );
  NAND2X2 U2496 ( .A(n2538), .B(n1987), .Y(n2389) );
  BUFX12 U2497 ( .A(n2343), .Y(n1975) );
  XNOR2X4 U2498 ( .A(n2024), .B(n1810), .Y(n2199) );
  NAND2BX2 U2499 ( .AN(\U4/temp7t[0] ), .B(\U4/U6/temp[0] ), .Y(n1455) );
  BUFX12 U2500 ( .A(n2405), .Y(n2560) );
  XOR2X4 U2501 ( .A(n2556), .B(n1725), .Y(n1722) );
  NAND2X4 U2502 ( .A(n1783), .B(n1790), .Y(n2311) );
  OAI2BB2X2 U2503 ( .B0(n2542), .B1(n1848), .A0N(n1848), .A1N(n2542), .Y(n2595) );
  CLKINVX3 U2504 ( .A(n2568), .Y(n812) );
  AOI2BB2X4 U2505 ( .B0(temp1t[3]), .B1(n1085), .A0N(n1085), .A1N(temp1t[3]), 
        .Y(n1846) );
  INVX8 U2506 ( .A(temp1t[4]), .Y(n1032) );
  XOR2X1 U2507 ( .A(n2787), .B(n2786), .Y(n2788) );
  OAI222X1 U2508 ( .A0(x0[2]), .A1(x7[2]), .B0(x0[2]), .B1(n572), .C0(x7[2]), 
        .C1(n572), .Y(n1223) );
  OAI222X1 U2509 ( .A0(x2[2]), .A1(x5[2]), .B0(x2[2]), .B1(n600), .C0(x5[2]), 
        .C1(n600), .Y(n1205) );
  XNOR3X2 U2510 ( .A(n2727), .B(\intadd_28/n1 ), .C(n2837), .Y(n2829) );
  NAND2X1 U2511 ( .A(n2732), .B(\intadd_28/n1 ), .Y(n2728) );
  NAND2X1 U2512 ( .A(n2809), .B(n2823), .Y(n2802) );
  XNOR3X2 U2513 ( .A(n2727), .B(n2749), .C(n2666), .Y(n2806) );
  XNOR3X2 U2514 ( .A(\U3/temp10t[8] ), .B(\U3/temp10t[7] ), .C(n2631), .Y(
        n2794) );
  NAND2BX1 U2515 ( .AN(\U3/temp10t[4] ), .B(\U3/temp10t[3] ), .Y(n2616) );
  OAI2BB1X4 U2516 ( .A0N(n2137), .A1N(n1310), .B0(n1008), .Y(n2340) );
  OAI21X2 U2517 ( .A0(n724), .A1(n852), .B0(n1520), .Y(n1266) );
  NAND2BX1 U2518 ( .AN(n2842), .B(n2770), .Y(n2767) );
  NAND2X1 U2519 ( .A(n2842), .B(n2783), .Y(n2406) );
  OAI2BB1X4 U2520 ( .A0N(n2692), .A1N(n2691), .B0(n2779), .Y(n2223) );
  NAND2X4 U2521 ( .A(n1664), .B(n743), .Y(n2452) );
  NAND2X4 U2522 ( .A(n1698), .B(n2565), .Y(n2421) );
  XNOR2X2 U2523 ( .A(n2266), .B(n2267), .Y(n1464) );
  INVX4 U2524 ( .A(n1467), .Y(n966) );
  NAND2X4 U2525 ( .A(n2494), .B(n659), .Y(n2306) );
  NAND2X4 U2526 ( .A(n660), .B(n1910), .Y(n2179) );
  NAND2X2 U2527 ( .A(n1917), .B(n1923), .Y(n2242) );
  OAI2BB1X4 U2528 ( .A0N(n992), .A1N(n1362), .B0(n996), .Y(n2310) );
  INVX8 U2529 ( .A(n1379), .Y(n996) );
  NAND2X4 U2530 ( .A(n637), .B(n1980), .Y(n2187) );
  NAND2X2 U2531 ( .A(n2579), .B(n1980), .Y(n2189) );
  INVX4 U2532 ( .A(n1978), .Y(n2345) );
  INVX4 U2533 ( .A(n2333), .Y(n2366) );
  OAI2BB1X4 U2534 ( .A0N(n743), .A1N(n736), .B0(n2446), .Y(n2445) );
  NAND2X4 U2535 ( .A(n1676), .B(n2561), .Y(n2173) );
  INVX8 U2536 ( .A(n2219), .Y(n2526) );
  XOR2X2 U2537 ( .A(n1767), .B(n1785), .Y(n2427) );
  AOI22X2 U2538 ( .A0(n1035), .A1(temp3t[5]), .B0(temp2t[5]), .B1(n1038), .Y(
        n1819) );
  XOR2X2 U2539 ( .A(n1797), .B(n1796), .Y(n2304) );
  NAND2X1 U2540 ( .A(n1085), .B(temp1t[3]), .Y(n2169) );
  INVX1 U2541 ( .A(temp3t[6]), .Y(n2278) );
  XOR2X1 U2542 ( .A(n2841), .B(n2790), .Y(n2791) );
  XOR2X1 U2543 ( .A(n2232), .B(n2839), .Y(n2819) );
  NAND2X1 U2544 ( .A(\intadd_28/n1 ), .B(n2752), .Y(n2746) );
  NAND2X1 U2545 ( .A(n2824), .B(n2823), .Y(n2828) );
  NAND2X2 U2546 ( .A(n2725), .B(n2644), .Y(n2645) );
  INVX1 U2547 ( .A(n2708), .Y(n2657) );
  NAND2X1 U2548 ( .A(n2795), .B(n2794), .Y(n2654) );
  NAND2BX1 U2549 ( .AN(\U3/temp10t[4] ), .B(\U3/temp10t[5] ), .Y(n2617) );
  NAND2BX1 U2550 ( .AN(\U3/temp10t[5] ), .B(\U3/temp10t[4] ), .Y(n2618) );
  OAI22X2 U2551 ( .A0(n691), .A1(n1513), .B0(n690), .B1(n1515), .Y(n1516) );
  AOI222X4 U2552 ( .A0(n690), .A1(n691), .B0(n690), .B1(n679), .C0(n691), .C1(
        n679), .Y(\U3/temp10[12] ) );
  MXI2X4 U2553 ( .A(n2476), .B(n2475), .S0(n2171), .Y(n2477) );
  XOR2X1 U2554 ( .A(n2775), .B(n2774), .Y(n2790) );
  XOR2X1 U2555 ( .A(n2770), .B(n2842), .Y(n2247) );
  OAI21X4 U2556 ( .A0(n2694), .A1(n2688), .B0(n2214), .Y(n2213) );
  XNOR3X2 U2557 ( .A(\U3/temp9t[7] ), .B(n2606), .C(n2682), .Y(n2779) );
  NOR2X1 U2558 ( .A(\U3/temp9t[2] ), .B(n2144), .Y(n2194) );
  NOR2X2 U2559 ( .A(\U3/temp11[1] ), .B(\U3/temp9t[1] ), .Y(n2193) );
  NAND2X4 U2560 ( .A(n1700), .B(n1638), .Y(n2391) );
  NAND2X4 U2561 ( .A(n1700), .B(n2557), .Y(n2390) );
  XOR2X4 U2562 ( .A(n1856), .B(n2494), .Y(n2502) );
  OAI21X1 U2563 ( .A0(n1493), .A1(\U4/U5/temp[6] ), .B0(n1019), .Y(n2268) );
  NAND2X4 U2564 ( .A(n654), .B(n2522), .Y(n2347) );
  NAND2X4 U2565 ( .A(n1868), .B(n659), .Y(n2307) );
  NAND2X4 U2566 ( .A(n2494), .B(n1868), .Y(n2305) );
  NAND2X2 U2567 ( .A(n2134), .B(n1874), .Y(n2203) );
  NAND2X2 U2568 ( .A(n2134), .B(n1875), .Y(n2204) );
  NAND2X2 U2569 ( .A(n1875), .B(n1874), .Y(n2205) );
  NAND2X4 U2570 ( .A(n660), .B(n2550), .Y(n2178) );
  NAND2X4 U2571 ( .A(n1893), .B(n752), .Y(n1890) );
  BUFX12 U2572 ( .A(n1885), .Y(n2550) );
  BUFX16 U2573 ( .A(n1942), .Y(n2589) );
  XOR2X4 U2574 ( .A(n2514), .B(n2520), .Y(\U1/temp_xxx[10] ) );
  INVX8 U2575 ( .A(n1981), .Y(n637) );
  OAI2BB2X4 U2576 ( .B0(n1994), .B1(n667), .A0N(n667), .A1N(n1994), .Y(n1972)
         );
  XOR2X2 U2577 ( .A(n2532), .B(n2007), .Y(n2005) );
  XOR2X4 U2578 ( .A(n2036), .B(n1948), .Y(n1989) );
  XOR2X4 U2579 ( .A(n1946), .B(n2037), .Y(n1997) );
  XOR2X4 U2580 ( .A(n2045), .B(n1851), .Y(n1951) );
  OAI2BB1X4 U2581 ( .A0N(n980), .A1N(n976), .B0(n2424), .Y(n2423) );
  XNOR2X2 U2582 ( .A(n1441), .B(n1452), .Y(n1415) );
  NAND2X4 U2583 ( .A(n737), .B(n1658), .Y(n2442) );
  INVX8 U2584 ( .A(n1683), .Y(n735) );
  NAND2X4 U2585 ( .A(n1755), .B(n2562), .Y(n2399) );
  NAND2X4 U2586 ( .A(n2556), .B(n1755), .Y(n2398) );
  XOR2X4 U2587 ( .A(n2586), .B(n2212), .Y(n1825) );
  XNOR2X4 U2588 ( .A(n2588), .B(n2548), .Y(n1773) );
  INVX8 U2589 ( .A(n2542), .Y(n2603) );
  OAI2BB1X4 U2590 ( .A0N(n800), .A1N(n2541), .B0(n787), .Y(n2570) );
  INVX1 U2591 ( .A(n1033), .Y(n2323) );
  NAND2BX1 U2592 ( .AN(n1032), .B(n1040), .Y(n2250) );
  CLKINVX3 U2593 ( .A(temp4t[4]), .Y(n1040) );
  XOR2X1 U2594 ( .A(n2714), .B(n2736), .Y(\U3/Ytt[1] ) );
  XOR2X1 U2595 ( .A(n2756), .B(n2755), .Y(n2757) );
  AOI222X4 U2596 ( .A0(x3[7]), .A1(x4[7]), .B0(x3[7]), .B1(n606), .C0(x4[7]), 
        .C1(n606), .Y(n1191) );
  NAND2X4 U2597 ( .A(n2838), .B(n2829), .Y(n2833) );
  OAI2BB1X4 U2598 ( .A0N(n2646), .A1N(n2733), .B0(n2645), .Y(n2729) );
  XNOR3X2 U2599 ( .A(\U3/temp10t[9] ), .B(\U3/temp10t[8] ), .C(n2629), .Y(
        n2667) );
  NAND2BX1 U2600 ( .AN(\U3/temp10t[6] ), .B(\U3/temp10t[5] ), .Y(n2620) );
  XNOR2X1 U2601 ( .A(n2295), .B(n2233), .Y(n2172) );
  OAI2BB1X2 U2602 ( .A0N(n1358), .A1N(n987), .B0(n2454), .Y(n2453) );
  INVX1 U2603 ( .A(n2772), .Y(n2775) );
  XOR2X1 U2604 ( .A(n2202), .B(n2763), .Y(n2764) );
  NAND2X4 U2605 ( .A(n2698), .B(n2697), .Y(n2244) );
  NOR2X1 U2606 ( .A(\U3/temp9t[3] ), .B(n2144), .Y(n2195) );
  AOI22X2 U2607 ( .A0(n2259), .A1(n1709), .B0(n749), .B1(n2555), .Y(n2258) );
  NAND2X2 U2608 ( .A(n2401), .B(n2565), .Y(n2422) );
  AND2X4 U2609 ( .A(n1486), .B(n1487), .Y(n2285) );
  NAND2X4 U2610 ( .A(n2522), .B(n658), .Y(n2349) );
  NAND2X4 U2611 ( .A(n1896), .B(n671), .Y(n2236) );
  INVX8 U2612 ( .A(n1375), .Y(n997) );
  INVX8 U2613 ( .A(n1984), .Y(n638) );
  NOR2X4 U2614 ( .A(n2587), .B(n1998), .Y(n2598) );
  NOR2X4 U2615 ( .A(n1997), .B(n1998), .Y(n2597) );
  INVX8 U2616 ( .A(n2532), .Y(n663) );
  XOR2X4 U2617 ( .A(n2043), .B(n1848), .Y(n1954) );
  OAI2BB1X2 U2618 ( .A0N(n980), .A1N(n1419), .B0(n984), .Y(n2471) );
  INVX8 U2619 ( .A(n1430), .Y(n981) );
  INVX8 U2620 ( .A(n1436), .Y(n984) );
  XNOR2X2 U2621 ( .A(n1453), .B(n1460), .Y(n1436) );
  INVX8 U2622 ( .A(n2529), .Y(n746) );
  OAI2BB1X4 U2623 ( .A0N(n2219), .A1N(n735), .B0(n2201), .Y(n2200) );
  INVX8 U2624 ( .A(n1684), .Y(n763) );
  INVX8 U2625 ( .A(n2146), .Y(n759) );
  XOR2X4 U2626 ( .A(n1825), .B(n1834), .Y(n1684) );
  NAND2X1 U2627 ( .A(n2548), .B(n2588), .Y(n2355) );
  INVX1 U2628 ( .A(n1808), .Y(n2342) );
  CLKBUFX8 U2629 ( .A(n766), .Y(n2576) );
  NAND2X1 U2630 ( .A(n1041), .B(temp1t[5]), .Y(n2281) );
  NAND2BX1 U2631 ( .AN(n1036), .B(n2278), .Y(n2277) );
  XOR2X1 U2632 ( .A(n2668), .B(n2825), .Y(\U3/Ytt[0] ) );
  XOR2X1 U2633 ( .A(n2817), .B(n2842), .Y(n2782) );
  NAND2X1 U2634 ( .A(n1237), .B(\U2/result1[3] ), .Y(n1259) );
  INVX1 U2635 ( .A(n2711), .Y(n2713) );
  INVX8 U2636 ( .A(\intadd_28/n1 ), .Y(n2823) );
  NAND2X2 U2637 ( .A(n2652), .B(n2725), .Y(n2649) );
  AOI2BB2X4 U2638 ( .B0(n2750), .B1(n2709), .A0N(n2729), .A1N(n2648), .Y(n2724) );
  OAI21X2 U2639 ( .A0(n2734), .A1(n2660), .B0(n2642), .Y(n2707) );
  NAND2BX1 U2640 ( .AN(\U3/temp10t[6] ), .B(\U3/temp10t[7] ), .Y(n2621) );
  NAND2BX1 U2641 ( .AN(\U3/temp10t[5] ), .B(\U3/temp10t[6] ), .Y(n2619) );
  NAND2BX1 U2642 ( .AN(\U3/temp10t[7] ), .B(\U3/temp10t[6] ), .Y(n2622) );
  OAI2BB1X4 U2643 ( .A0N(n1302), .A1N(n1315), .B0(n2272), .Y(n2271) );
  OAI21X4 U2644 ( .A0(n1302), .A1(n1315), .B0(n2273), .Y(n2272) );
  INVX8 U2645 ( .A(n1318), .Y(n1003) );
  INVX8 U2646 ( .A(n1321), .Y(n1005) );
  AFHCONX4 U2647 ( .A(n2841), .B(n2790), .CI(n2792), .CON(n2789) );
  INVX1 U2648 ( .A(n2687), .Y(n2693) );
  XOR2X1 U2649 ( .A(n2813), .B(n2812), .Y(n2814) );
  NOR2X1 U2650 ( .A(\U3/temp9t[4] ), .B(n2144), .Y(n2672) );
  AOI2BB2X4 U2651 ( .B0(n2534), .B1(n2510), .A0N(n2131), .A1N(n2511), .Y(n2509) );
  NAND2X4 U2652 ( .A(n2523), .B(n743), .Y(n2451) );
  NAND2X4 U2653 ( .A(n2523), .B(n1664), .Y(n2450) );
  NAND2X2 U2654 ( .A(n1638), .B(n2557), .Y(n2392) );
  OAI21X4 U2655 ( .A0(n731), .A1(n1703), .B0(n1702), .Y(n2356) );
  AOI2BB2X1 U2656 ( .B0(n1729), .B1(n2561), .A0N(n1729), .A1N(n2561), .Y(n1707) );
  AND2X4 U2657 ( .A(n1486), .B(n973), .Y(n2284) );
  NAND3X4 U2658 ( .A(n2305), .B(n2306), .C(n2307), .Y(n2308) );
  NAND2X2 U2659 ( .A(n2547), .B(n652), .Y(n2262) );
  AOI2BB2X4 U2660 ( .B0(n1905), .B1(n668), .A0N(n1905), .A1N(n668), .Y(n1859)
         );
  AND2X4 U2661 ( .A(n2130), .B(n1903), .Y(n2329) );
  NAND2X4 U2662 ( .A(n1897), .B(n1896), .Y(n2235) );
  XOR2X4 U2663 ( .A(n1917), .B(n1918), .Y(n1896) );
  NAND2X4 U2664 ( .A(n1961), .B(n640), .Y(n2491) );
  NAND2X4 U2665 ( .A(n1965), .B(n1957), .Y(n2464) );
  NAND2X4 U2666 ( .A(n1973), .B(n2380), .Y(n2429) );
  NAND2X4 U2667 ( .A(n1975), .B(n2538), .Y(n2388) );
  XOR2X4 U2668 ( .A(n2161), .B(n2011), .Y(n2008) );
  NAND2X4 U2669 ( .A(n1975), .B(n1987), .Y(n2387) );
  AOI2BB2X4 U2670 ( .B0(n2344), .B1(n1977), .A0N(n2346), .A1N(n2345), .Y(n2343) );
  XOR2X4 U2671 ( .A(n667), .B(n2000), .Y(n1999) );
  NAND2X4 U2672 ( .A(n2127), .B(n667), .Y(n2324) );
  NAND2X4 U2673 ( .A(n752), .B(n676), .Y(n1993) );
  XOR2X4 U2674 ( .A(n1949), .B(n2040), .Y(n2016) );
  OAI21X4 U2675 ( .A0(n2569), .A1(n1953), .B0(n2042), .Y(n2037) );
  INVX8 U2676 ( .A(n1427), .Y(n979) );
  XOR2X4 U2677 ( .A(n1719), .B(n2434), .Y(n2405) );
  AOI2BB2X4 U2678 ( .B0(n1739), .B1(n2537), .A0N(n1739), .A1N(n2537), .Y(n1670) );
  OAI2BB1X4 U2679 ( .A0N(n761), .A1N(n1771), .B0(n2132), .Y(n2218) );
  INVX8 U2680 ( .A(n1240), .Y(n764) );
  INVX8 U2681 ( .A(n1838), .Y(n766) );
  XOR2X4 U2682 ( .A(n1810), .B(n1811), .Y(n1784) );
  XOR2X1 U2683 ( .A(n2710), .B(n2713), .Y(n2668) );
  XOR2X1 U2684 ( .A(n2806), .B(\intadd_28/n1 ), .Y(n2807) );
  NAND2X1 U2685 ( .A(n574), .B(x7[0]), .Y(n1140) );
  NAND2X1 U2686 ( .A(n602), .B(x5[0]), .Y(n1172) );
  AOI222X1 U2687 ( .A0(x4[7]), .A1(n604), .B0(x4[7]), .B1(n1176), .C0(n604), 
        .C1(n1176), .Y(n1174) );
  AOI222X1 U2688 ( .A0(x6[7]), .A1(n576), .B0(x6[7]), .B1(n1144), .C0(n576), 
        .C1(n1144), .Y(n1142) );
  NAND2X4 U2689 ( .A(n2831), .B(n2830), .Y(n2832) );
  AOI2BB2X4 U2690 ( .B0(n2830), .B1(n2739), .A0N(n2738), .A1N(n2737), .Y(n2762) );
  OAI2BB1X2 U2691 ( .A0N(n2711), .A1N(n2824), .B0(n2710), .Y(n2712) );
  AOI2BB2X4 U2692 ( .B0(n2667), .B1(n2750), .A0N(n2748), .A1N(n2651), .Y(n2793) );
  OAI2BB1X4 U2693 ( .A0N(n2650), .A1N(n2724), .B0(n2649), .Y(n2748) );
  NAND2BX1 U2694 ( .AN(\U3/temp10t[9] ), .B(\U3/temp11[0] ), .Y(n2627) );
  NAND2BX1 U2695 ( .AN(\U3/temp10t[8] ), .B(\U3/temp10t[9] ), .Y(n2625) );
  NAND2BX1 U2696 ( .AN(\U3/temp10t[7] ), .B(\U3/temp10t[8] ), .Y(n2623) );
  INVX1 U2697 ( .A(\U3/temp10t[1] ), .Y(n2608) );
  NAND2BX1 U2698 ( .AN(\U3/temp10t[8] ), .B(\U3/temp10t[7] ), .Y(n2624) );
  NAND2BX1 U2699 ( .AN(\U3/temp10t[9] ), .B(\U3/temp10t[8] ), .Y(n2626) );
  NAND2BX1 U2700 ( .AN(\U3/temp11[0] ), .B(\U3/temp10t[9] ), .Y(n2628) );
  XOR2X1 U2701 ( .A(n1405), .B(\intadd_41/n1 ), .Y(\U4/temp7[10] ) );
  BUFX12 U2702 ( .A(n2271), .Y(n1313) );
  INVX8 U2703 ( .A(\intadd_35/n1 ), .Y(n679) );
  OAI21X1 U2704 ( .A0(n2551), .A1(n852), .B0(\U5/temp1[0] ), .Y(n1518) );
  INVX8 U2705 ( .A(\U5/temp2[0] ), .Y(n852) );
  XNOR2X4 U2706 ( .A(n2525), .B(n2499), .Y(n2485) );
  NAND2BX4 U2707 ( .AN(n2698), .B(n2780), .Y(n2245) );
  NOR2X4 U2708 ( .A(n2781), .B(n2779), .Y(n2225) );
  AOI2BB2X4 U2709 ( .B0(n2220), .B1(n2142), .A0N(n2213), .A1N(n2689), .Y(n2772) );
  NOR2X1 U2710 ( .A(\U3/temp9t[7] ), .B(n2144), .Y(n2675) );
  NOR2X1 U2711 ( .A(\U3/temp9t[6] ), .B(n2144), .Y(n2674) );
  NOR2X1 U2712 ( .A(\U3/temp9t[5] ), .B(n2144), .Y(n2673) );
  NAND2X4 U2713 ( .A(n2123), .B(n2558), .Y(n2460) );
  NAND2X4 U2714 ( .A(n2123), .B(n727), .Y(n2459) );
  AND2X4 U2715 ( .A(n728), .B(n744), .Y(n2433) );
  OAI21X4 U2716 ( .A0(n728), .A1(n744), .B0(n2524), .Y(n2432) );
  OAI21XL U2717 ( .A0(n752), .A1(n2566), .B0(n1730), .Y(n1817) );
  NAND2X4 U2718 ( .A(n967), .B(n965), .Y(n2318) );
  NAND2X4 U2719 ( .A(n967), .B(n1480), .Y(n2319) );
  OAI2BB1X4 U2720 ( .A0N(n1467), .A1N(n969), .B0(n2289), .Y(n2288) );
  OAI21X4 U2721 ( .A0(\U4/temp5t[0] ), .A1(\U4/U5/temp[0] ), .B0(n970), .Y(
        n1509) );
  INVX8 U2722 ( .A(n2495), .Y(n1882) );
  OAI2BB2X4 U2723 ( .B0(n1853), .B1(n2494), .A0N(n1856), .A1N(n2493), .Y(n2495) );
  OAI2BB2X4 U2724 ( .B0(n2547), .B1(n2482), .A0N(n2533), .A1N(n2481), .Y(n2483) );
  BUFX12 U2725 ( .A(n1865), .Y(n2552) );
  XOR2X4 U2726 ( .A(n668), .B(n1904), .Y(n1902) );
  AND2X4 U2727 ( .A(n1897), .B(n671), .Y(n2237) );
  NAND2X4 U2728 ( .A(n1961), .B(n643), .Y(n2490) );
  NAND2BX2 U2729 ( .AN(n989), .B(n2249), .Y(n2248) );
  XOR2X4 U2730 ( .A(n1961), .B(n2538), .Y(n2488) );
  NAND2X4 U2731 ( .A(n1965), .B(n2346), .Y(n2465) );
  NAND2X4 U2732 ( .A(n1968), .B(n1966), .Y(n2437) );
  NAND2X4 U2733 ( .A(n1968), .B(n1969), .Y(n2438) );
  NAND2X4 U2734 ( .A(n1973), .B(n646), .Y(n2430) );
  NOR2X4 U2735 ( .A(n639), .B(n2031), .Y(n1984) );
  XOR2X2 U2736 ( .A(n1989), .B(n1990), .Y(n1988) );
  OR2X4 U2737 ( .A(n2127), .B(n667), .Y(n2326) );
  XOR2X4 U2738 ( .A(n2033), .B(n1939), .Y(n2015) );
  NAND2X4 U2739 ( .A(n2026), .B(n833), .Y(n2215) );
  BUFX16 U2740 ( .A(n1285), .Y(n2567) );
  AOI22X2 U2741 ( .A0(n2138), .A1(n1414), .B0(n975), .B1(n1415), .Y(n1413) );
  OAI2BB1X2 U2742 ( .A0N(n1415), .A1N(n981), .B0(n2361), .Y(n2360) );
  NAND2X4 U2743 ( .A(n1751), .B(n1715), .Y(n2402) );
  OAI2BB1X4 U2744 ( .A0N(n2545), .A1N(n2129), .B0(n2505), .Y(n2504) );
  INVX8 U2745 ( .A(n1653), .Y(n736) );
  INVX8 U2746 ( .A(n1657), .Y(n737) );
  NAND2X4 U2747 ( .A(n1685), .B(n747), .Y(n1661) );
  INVX8 U2748 ( .A(n2557), .Y(n747) );
  BUFX12 U2749 ( .A(n1686), .Y(n2557) );
  AOI22X4 U2750 ( .A0(n2156), .A1(n2369), .B0(n1744), .B1(n2219), .Y(n2368) );
  AOI22X4 U2751 ( .A0(n2561), .A1(n2228), .B0(n1730), .B1(n748), .Y(n1735) );
  XOR2X4 U2752 ( .A(n1777), .B(n2358), .Y(n1775) );
  XOR2X4 U2753 ( .A(n2414), .B(n2135), .Y(n1724) );
  OAI2BB1X4 U2754 ( .A0N(n2124), .A1N(n1834), .B0(n2287), .Y(n2286) );
  NAND2X2 U2755 ( .A(n2586), .B(n2124), .Y(n2287) );
  NAND2X4 U2756 ( .A(n764), .B(n1955), .Y(n1828) );
  INVX8 U2757 ( .A(n2601), .Y(n1955) );
  INVX8 U2758 ( .A(n1850), .Y(n1123) );
  AOI2BB2X4 U2759 ( .B0(temp2t[2]), .B1(temp3t[2]), .A0N(temp3t[2]), .A1N(
        temp2t[2]), .Y(n1851) );
  XNOR2X1 U2760 ( .A(n2842), .B(n2783), .Y(n2784) );
  XOR2X1 U2761 ( .A(n2824), .B(n2823), .Y(n2805) );
  NAND2X2 U2762 ( .A(n2760), .B(n2759), .Y(n2742) );
  OAI2BB1X4 U2763 ( .A0N(n2654), .A1N(n2793), .B0(n2653), .Y(n2666) );
  NAND2X2 U2764 ( .A(n2703), .B(n2652), .Y(n2653) );
  NAND2BX1 U2765 ( .AN(\U3/temp11[0] ), .B(\U3/temp11[1] ), .Y(n2662) );
  OAI2BB1X4 U2766 ( .A0N(n2639), .A1N(n2610), .B0(n2609), .Y(n2641) );
  NAND2BX1 U2767 ( .AN(\U3/temp11[1] ), .B(\U3/temp11[0] ), .Y(n2664) );
  NAND2BX1 U2768 ( .AN(n1002), .B(n2137), .Y(n2457) );
  OAI2BB1X4 U2769 ( .A0N(n2425), .A1N(n2170), .B0(n2426), .Y(n2171) );
  NAND2BX4 U2770 ( .AN(\U5/temp7t[0] ), .B(\U5/U6/temp[0] ), .Y(n1346) );
  NAND2X4 U2771 ( .A(n2816), .B(n2839), .Y(n2415) );
  OAI21XL U2772 ( .A0(n2670), .A1(n2689), .B0(n2693), .Y(n2234) );
  CLKINVX3 U2773 ( .A(n2778), .Y(n2786) );
  NAND2X2 U2774 ( .A(n2763), .B(n2773), .Y(n2222) );
  XOR2X1 U2775 ( .A(n2686), .B(n2685), .Y(n2694) );
  NOR2X1 U2776 ( .A(\U3/temp12[1] ), .B(n2144), .Y(n2695) );
  NOR2X1 U2777 ( .A(\U3/temp12[0] ), .B(n2144), .Y(n2678) );
  NOR2X1 U2778 ( .A(\U3/temp9t[9] ), .B(n2144), .Y(n2677) );
  NOR2X1 U2779 ( .A(\U3/temp9t[8] ), .B(n2144), .Y(n2676) );
  NAND2X2 U2780 ( .A(n727), .B(n2558), .Y(n2461) );
  OAI2BB1X4 U2781 ( .A0N(n1463), .A1N(n1469), .B0(n973), .Y(n2467) );
  OAI2BB1X4 U2782 ( .A0N(n968), .A1N(n1471), .B0(n2141), .Y(n2463) );
  BUFX12 U2783 ( .A(n2410), .Y(n1474) );
  OAI2BB1X4 U2784 ( .A0N(n1463), .A1N(n1476), .B0(n2411), .Y(n2410) );
  OAI2BB1X4 U2785 ( .A0N(n968), .A1N(n964), .B0(n2412), .Y(n2411) );
  INVX8 U2786 ( .A(n2483), .Y(n1856) );
  OAI21X4 U2787 ( .A0(n1906), .A1(n2540), .B0(n1909), .Y(n2274) );
  NAND2X4 U2788 ( .A(n1906), .B(n2540), .Y(n2275) );
  NAND3BX4 U2789 ( .AN(n2237), .B(n2235), .C(n2236), .Y(n2238) );
  MX2X2 U2790 ( .A(n2594), .B(n760), .S0(n678), .Y(n2164) );
  BUFX12 U2791 ( .A(n1900), .Y(n2527) );
  AOI22X4 U2792 ( .A0(n1959), .A1(n2515), .B0(n1957), .B1(n2536), .Y(n2514) );
  CLKINVX3 U2793 ( .A(n1373), .Y(n993) );
  XNOR2X2 U2794 ( .A(n1387), .B(n1388), .Y(n1375) );
  NAND2BX4 U2795 ( .AN(\U5/temp5t[0] ), .B(\U5/U5/temp[0] ), .Y(n1398) );
  AOI2BB2X4 U2796 ( .B0(n2008), .B1(n2333), .A0N(n2008), .A1N(n2333), .Y(n1962) );
  OAI2BB2X4 U2797 ( .B0(n1999), .B1(n664), .A0N(n1999), .A1N(n664), .Y(n1964)
         );
  OAI2BB1X4 U2798 ( .A0N(n2161), .A1N(n2011), .B0(n2366), .Y(n2365) );
  NOR2X4 U2799 ( .A(n666), .B(n2532), .Y(n2270) );
  AOI21X4 U2800 ( .A0(n666), .A1(n2532), .B0(n2007), .Y(n2269) );
  OR3X4 U2801 ( .A(n2596), .B(n2597), .C(n2598), .Y(n1990) );
  XOR2X2 U2802 ( .A(n1953), .B(n1954), .Y(n1944) );
  INVX8 U2803 ( .A(n2016), .Y(n2587) );
  XOR2X4 U2804 ( .A(n1926), .B(n1930), .Y(n1914) );
  XNOR2X4 U2805 ( .A(n665), .B(n1922), .Y(n2333) );
  XNOR2X4 U2806 ( .A(n2023), .B(n1798), .Y(n1923) );
  NAND2X4 U2807 ( .A(n2018), .B(n1930), .Y(n2230) );
  NAND2X4 U2808 ( .A(n2018), .B(n1926), .Y(n2229) );
  NAND2X4 U2809 ( .A(n2026), .B(n1928), .Y(n2216) );
  MXI2X4 U2810 ( .A(n724), .B(n2567), .S0(n1123), .Y(n1953) );
  INVX4 U2811 ( .A(n2567), .Y(n724) );
  XNOR2X4 U2812 ( .A(n2044), .B(n1852), .Y(n1952) );
  INVX8 U2813 ( .A(n1414), .Y(n975) );
  OAI21X4 U2814 ( .A0(n980), .A1(n1419), .B0(n2471), .Y(n2470) );
  CLKINVX3 U2815 ( .A(n1424), .Y(n976) );
  OAI2BB1X4 U2816 ( .A0N(n2138), .A1N(n2359), .B0(n2360), .Y(n1427) );
  CLKINVX3 U2817 ( .A(n981), .Y(n2359) );
  MXI2X4 U2818 ( .A(n726), .B(n739), .S0(n728), .Y(n2507) );
  CLKINVX3 U2819 ( .A(n2565), .Y(n2314) );
  NAND2X2 U2820 ( .A(n2126), .B(n2556), .Y(n2386) );
  INVX8 U2821 ( .A(n1770), .Y(n733) );
  NOR2X4 U2822 ( .A(n752), .B(n1687), .Y(n1680) );
  MXI2X4 U2823 ( .A(n2584), .B(n1826), .S0(n1827), .Y(n1687) );
  NAND2X2 U2824 ( .A(n2556), .B(n2562), .Y(n2397) );
  NAND2X4 U2825 ( .A(n1783), .B(n2528), .Y(n2312) );
  NAND2X4 U2826 ( .A(n1778), .B(n1780), .Y(n2377) );
  NAND2X4 U2827 ( .A(n1778), .B(n2159), .Y(n2376) );
  OR2X4 U2828 ( .A(n2575), .B(n768), .Y(n2335) );
  AOI21X4 U2829 ( .A0(n2575), .A1(n768), .B0(n2574), .Y(n2334) );
  INVX8 U2830 ( .A(n1805), .Y(n2575) );
  AOI2BB2X4 U2831 ( .B0(n2564), .B1(n2190), .A0N(n2191), .A1N(n2192), .Y(n1832) );
  INVX8 U2832 ( .A(n2559), .Y(n775) );
  XOR2X4 U2833 ( .A(n1852), .B(n1847), .Y(n1838) );
  CLKBUFX8 U2834 ( .A(n1839), .Y(n2559) );
  AOI22X2 U2835 ( .A0(n1850), .A1(n2551), .B0(n787), .B1(n1123), .Y(n1839) );
  AOI2BB2X4 U2836 ( .B0(temp1t[1]), .B1(temp4t[1]), .A0N(temp4t[1]), .A1N(
        temp1t[1]), .Y(n1850) );
  AOI22X4 U2837 ( .A0(temp2t[3]), .A1(n1083), .B0(temp3t[3]), .B1(n1081), .Y(
        n1844) );
  NAND2X1 U2838 ( .A(n962), .B(temp1t[7]), .Y(n2371) );
  NAND2BX1 U2839 ( .AN(temp4t[6]), .B(n2323), .Y(n2322) );
  NAND2X4 U2840 ( .A(n1843), .B(n1085), .Y(n2168) );
  NAND2X4 U2841 ( .A(n1841), .B(n1083), .Y(n2208) );
  NAND2X4 U2842 ( .A(n1845), .B(n1080), .Y(n2197) );
  NAND2X4 U2843 ( .A(n1845), .B(temp3t[2]), .Y(n2196) );
  INVX1 U2844 ( .A(\intadd_38/SUM[4] ), .Y(n794) );
  INVX1 U2845 ( .A(\intadd_41/SUM[4] ), .Y(n817) );
  XOR2X1 U2846 ( .A(\intadd_28/n1 ), .B(n2752), .Y(n2753) );
  XOR2X1 U2847 ( .A(\intadd_28/n1 ), .B(n2796), .Y(n2751) );
  XOR2X4 U2848 ( .A(n2835), .B(n2834), .Y(n2844) );
  MXI2X4 U2849 ( .A(n2833), .B(n2832), .S0(\intadd_28/n1 ), .Y(n2835) );
  AOI2BB2X4 U2850 ( .B0(n2823), .B1(n2799), .A0N(n2798), .A1N(n2797), .Y(n2810) );
  XNOR3X4 U2851 ( .A(\intadd_28/n1 ), .B(n2732), .C(n2731), .Y(n2760) );
  AOI2BB2X4 U2852 ( .B0(n2823), .B1(n2727), .A0N(n2837), .A1N(n2726), .Y(n2731) );
  NAND2BX1 U2853 ( .AN(\U3/temp11[1] ), .B(n2144), .Y(n2699) );
  NAND2X1 U2854 ( .A(\U3/temp11[1] ), .B(n2606), .Y(n2701) );
  AOI2BB2X4 U2855 ( .B0(n2727), .B1(n2667), .A0N(n2666), .A1N(n2665), .Y(n2705) );
  OAI2BB1X4 U2856 ( .A0N(n2618), .A1N(n2634), .B0(n2617), .Y(n2633) );
  OAI2BB1X4 U2857 ( .A0N(n2616), .A1N(n2636), .B0(n2615), .Y(n2634) );
  OAI2BB1X4 U2858 ( .A0N(n2614), .A1N(n2637), .B0(n2613), .Y(n2636) );
  OAI2BB1X4 U2859 ( .A0N(n2612), .A1N(n2641), .B0(n2611), .Y(n2637) );
  OAI21X4 U2860 ( .A0(n2137), .A1(n1310), .B0(n2340), .Y(n1308) );
  OAI21X2 U2861 ( .A0(\U5/temp7t[0] ), .A1(\U5/U6/temp[0] ), .B0(n1006), .Y(
        n1348) );
  INVX8 U2862 ( .A(n1517), .Y(n785) );
  MXI2X4 U2863 ( .A(n2500), .B(n2501), .S0(n2592), .Y(\U1/temp_xxx[9] ) );
  AOI2BB2X4 U2864 ( .B0(n2719), .B1(n2136), .A0N(n2718), .A1N(n2296), .Y(n2295) );
  OAI2BB1X4 U2865 ( .A0N(n2244), .A1N(n2766), .B0(n2245), .Y(n2718) );
  AOI2BB2X4 U2866 ( .B0(n2779), .B1(n2781), .A0N(n2225), .A1N(n2697), .Y(n2811) );
  OAI2BB1X4 U2867 ( .A0N(n2769), .A1N(n2142), .B0(n2223), .Y(n2765) );
  INVX8 U2868 ( .A(n2691), .Y(n2769) );
  OAI2BB1X4 U2869 ( .A0N(n2221), .A1N(n2772), .B0(n2222), .Y(n2691) );
  INVX8 U2870 ( .A(n2210), .Y(n2763) );
  INVX8 U2871 ( .A(n2202), .Y(n2812) );
  NAND2X2 U2872 ( .A(n2813), .B(n2202), .Y(n2226) );
  AOI2BB2X4 U2873 ( .B0(\U3/temp11[1] ), .B1(\U3/temp9t[1] ), .A0N(n2193), 
        .A1N(n2669), .Y(n2686) );
  OAI2BB1X2 U2874 ( .A0N(n2133), .A1N(n1664), .B0(n739), .Y(n2511) );
  CLKINVX3 U2875 ( .A(n2512), .Y(n2513) );
  OAI2BB1X2 U2876 ( .A0N(n738), .A1N(n1664), .B0(n2530), .Y(n2512) );
  AND3X4 U2877 ( .A(n2339), .B(n2338), .C(n2337), .Y(n1702) );
  CLKINVX3 U2878 ( .A(n2517), .Y(n2518) );
  OR2X4 U2879 ( .A(n1469), .B(n1463), .Y(n2468) );
  BUFX12 U2880 ( .A(n2462), .Y(n1469) );
  AOI2BB2X4 U2881 ( .B0(n2535), .B1(n2447), .A0N(n1853), .A1N(n2134), .Y(n2533) );
  BUFX12 U2882 ( .A(n1862), .Y(n2549) );
  CLKINVX3 U2883 ( .A(n1853), .Y(n2482) );
  NAND3BX4 U2884 ( .AN(n2329), .B(n2327), .C(n2328), .Y(n2330) );
  CLKINVX3 U2885 ( .A(n1947), .Y(n2572) );
  CLKINVX3 U2886 ( .A(n1949), .Y(n2593) );
  XOR2X4 U2887 ( .A(n1913), .B(n1914), .Y(n1910) );
  INVX8 U2888 ( .A(n2540), .Y(n670) );
  BUFX12 U2889 ( .A(n1899), .Y(n2540) );
  AOI222X4 U2890 ( .A0(n1951), .A1(n1952), .B0(n1951), .B1(n1945), .C0(n1945), 
        .C1(n1952), .Y(n1947) );
  INVX8 U2891 ( .A(n2456), .Y(n1352) );
  OAI2BB2X4 U2892 ( .B0(n992), .B1(n1358), .A0N(n987), .A1N(n2455), .Y(n2456)
         );
  OAI22X4 U2893 ( .A0(n1360), .A1(n2428), .B0(n1354), .B1(n1375), .Y(n1357) );
  OAI21X4 U2894 ( .A0(n992), .A1(n1362), .B0(n2310), .Y(n1360) );
  AOI22X4 U2895 ( .A0(n991), .A1(n2248), .B0(n989), .B1(n1371), .Y(n1367) );
  OAI2BB1X4 U2896 ( .A0N(n2176), .A1N(n1373), .B0(n2177), .Y(n1370) );
  OAI21X2 U2897 ( .A0(\U5/temp5t[0] ), .A1(\U5/U5/temp[0] ), .B0(n994), .Y(
        n1400) );
  XOR2X4 U2898 ( .A(n2012), .B(n2379), .Y(n2413) );
  OAI222X4 U2899 ( .A0(n2002), .A1(n2004), .B0(n2002), .B1(n664), .C0(n2004), 
        .C1(n664), .Y(n2013) );
  BUFX12 U2900 ( .A(n2006), .Y(n2532) );
  NAND2X2 U2901 ( .A(n833), .B(n1928), .Y(n2217) );
  INVX8 U2902 ( .A(n2599), .Y(n1950) );
  XOR2X2 U2903 ( .A(n2046), .B(n2600), .Y(n2599) );
  AOI22X4 U2904 ( .A0(n975), .A1(n2503), .B0(n1411), .B1(n2138), .Y(n1409) );
  OAI21X4 U2905 ( .A0(n2470), .A1(n1411), .B0(n2489), .Y(n1414) );
  OAI2BB1X4 U2906 ( .A0N(n1424), .A1N(n1411), .B0(n2423), .Y(n1422) );
  CLKINVX3 U2907 ( .A(n739), .Y(n2505) );
  OAI2BB1X4 U2908 ( .A0N(n2443), .A1N(n2444), .B0(n2445), .Y(n1650) );
  CLKINVX3 U2909 ( .A(n736), .Y(n2444) );
  OAI2BB1X4 U2910 ( .A0N(n2314), .A1N(n2315), .B0(n2316), .Y(n1657) );
  CLKINVX3 U2911 ( .A(n746), .Y(n2315) );
  CLKINVX3 U2912 ( .A(n743), .Y(n2443) );
  XOR2X4 U2913 ( .A(n1754), .B(n2562), .Y(n1651) );
  AOI22X4 U2914 ( .A0(n2332), .A1(n733), .B0(n2553), .B1(n2157), .Y(n2331) );
  OAI2BB1X4 U2915 ( .A0N(n2526), .A1N(n1683), .B0(n2200), .Y(n1771) );
  INVX4 U2916 ( .A(n1744), .Y(n762) );
  XOR2X4 U2917 ( .A(n1713), .B(n1714), .Y(n1633) );
  XOR2X4 U2918 ( .A(n1772), .B(n1773), .Y(n1744) );
  XNOR2X4 U2919 ( .A(n1824), .B(n1825), .Y(n1673) );
  XOR2X2 U2920 ( .A(n1805), .B(n1837), .Y(n1737) );
  OAI21X2 U2921 ( .A0(n1240), .A1(n1955), .B0(n1826), .Y(n1688) );
  XNOR2X4 U2922 ( .A(n2159), .B(n1780), .Y(n1769) );
  BUFX12 U2923 ( .A(n1724), .Y(n2556) );
  OAI2BB2X4 U2924 ( .B0(n2293), .B1(n2162), .A0N(n1776), .A1N(n2292), .Y(n2294) );
  NAND2X2 U2925 ( .A(n2162), .B(n2293), .Y(n2292) );
  NAND2BX4 U2926 ( .AN(n2334), .B(n2335), .Y(n2336) );
  XNOR2X4 U2927 ( .A(n1786), .B(n1787), .Y(n1767) );
  INVX4 U2928 ( .A(n1807), .Y(n2582) );
  AOI22X4 U2929 ( .A0(temp1t[2]), .A1(temp4t[2]), .B0(n1084), .B1(n1079), .Y(
        n1852) );
  INVX8 U2930 ( .A(n2595), .Y(n1829) );
  OAI22X4 U2931 ( .A0(n1121), .A1(temp3t[1]), .B0(n1122), .B1(temp2t[1]), .Y(
        n1848) );
  AOI21X4 U2932 ( .A0(n812), .A1(n2602), .B0(n2603), .Y(n2601) );
  XOR2X2 U2933 ( .A(n1851), .B(n1845), .Y(n1833) );
  BUFX12 U2934 ( .A(n1784), .Y(n2528) );
  AOI2BB2X4 U2935 ( .B0(n1807), .B1(n2322), .A0N(n1042), .A1N(n2323), .Y(n2321) );
  NAND2X4 U2936 ( .A(n1843), .B(temp1t[3]), .Y(n2167) );
  NAND2X4 U2937 ( .A(n1820), .B(n1034), .Y(n2256) );
  NAND2X4 U2938 ( .A(n1820), .B(temp3t[4]), .Y(n2255) );
  NAND2X4 U2939 ( .A(n1841), .B(temp2t[3]), .Y(n2207) );
  NAND2X4 U2940 ( .A(n850), .B(n2568), .Y(n1849) );
  INVX1 U2941 ( .A(\U2/result1[11] ), .Y(n888) );
  AFHCONX2 U2942 ( .A(x6[8]), .B(n575), .CI(n1142), .CON(temp7[9]) );
  AFHCONX2 U2943 ( .A(x4[8]), .B(n603), .CI(n1174), .CON(temp5[9]) );
  AOI2BB2X4 U2944 ( .B0(n2823), .B1(n2804), .A0N(n2808), .A1N(n2803), .Y(n2827) );
  OAI2BB1X4 U2945 ( .A0N(n2802), .A1N(n2810), .B0(n2801), .Y(n2808) );
  AOI2BB2X4 U2946 ( .B0(n2745), .B1(n2744), .A0N(n2758), .A1N(n2743), .Y(n2754) );
  OAI2BB1X4 U2947 ( .A0N(n2742), .A1N(n2762), .B0(n2741), .Y(n2758) );
  CLKINVX3 U2948 ( .A(n2736), .Y(n2739) );
  OAI2BB1X4 U2949 ( .A0N(n2713), .A1N(n2825), .B0(n2712), .Y(n2736) );
  INVX8 U2950 ( .A(n2824), .Y(n2825) );
  OAI2BB1X4 U2951 ( .A0N(n2706), .A1N(n2705), .B0(n2704), .Y(n2837) );
  XNOR3X4 U2952 ( .A(n2702), .B(n2795), .C(n2705), .Y(n2824) );
  NAND2X2 U2953 ( .A(n2708), .B(n2655), .Y(n2660) );
  INVX1 U2954 ( .A(\U3/temp10t[2] ), .Y(n2638) );
  INVX1 U2955 ( .A(\U3/temp10t[4] ), .Y(n2635) );
  OAI2BB1X4 U2956 ( .A0N(n2626), .A1N(n2629), .B0(n2625), .Y(n2630) );
  OAI2BB1X4 U2957 ( .A0N(n2624), .A1N(n2631), .B0(n2623), .Y(n2629) );
  OAI2BB1X4 U2958 ( .A0N(n2622), .A1N(n2632), .B0(n2621), .Y(n2631) );
  OAI2BB1X4 U2959 ( .A0N(n2620), .A1N(n2633), .B0(n2619), .Y(n2632) );
  AOI21X1 U2960 ( .A0(n1252), .A1(n931), .B0(n1233), .Y(\intadd_44/B[3] ) );
  INVX8 U2961 ( .A(n1305), .Y(n999) );
  OAI21X4 U2962 ( .A0(n1308), .A1(n2448), .B0(n2449), .Y(n1305) );
  AOI21X4 U2963 ( .A0(\U5/temp7t[0] ), .A1(\U5/U6/temp[0] ), .B0(n1348), .Y(
        n1337) );
  XOR2X2 U2964 ( .A(n1349), .B(n1350), .Y(n1312) );
  AOI222X4 U2965 ( .A0(\U5/temp1[1] ), .A1(n1099), .B0(n1281), .B1(
        \U5/temp1[1] ), .C0(n1099), .C1(n1281), .Y(n1517) );
  AOI2BB2X4 U2966 ( .B0(n2232), .B1(n2842), .A0N(n2820), .A1N(n2419), .Y(n2170) );
  OAI2BB1X4 U2967 ( .A0N(n2417), .A1N(n2822), .B0(n2418), .Y(n2820) );
  NAND2BX4 U2968 ( .AN(n2234), .B(n2232), .Y(n2722) );
  XOR2X4 U2969 ( .A(n2771), .B(n2247), .Y(n2841) );
  XNOR3X4 U2970 ( .A(n2233), .B(n2780), .C(n2698), .Y(n2232) );
  INVX4 U2971 ( .A(n2697), .Y(n2780) );
  OAI2BB1X4 U2972 ( .A0N(n2226), .A1N(n2811), .B0(n2227), .Y(n2698) );
  AOI2BB2X4 U2973 ( .B0(n2812), .B1(n2763), .A0N(n2765), .A1N(n2224), .Y(n2781) );
  INVX1 U2974 ( .A(\U3/temp9t[6] ), .Y(n2211) );
  INVX8 U2975 ( .A(n2842), .Y(n2839) );
  AOI2BB2X4 U2976 ( .B0(n2144), .B1(\U3/temp9t[9] ), .A0N(n2679), .A1N(n2677), 
        .Y(n2680) );
  AOI2BB2X4 U2977 ( .B0(n2144), .B1(\U3/temp9t[7] ), .A0N(n2682), .A1N(n2675), 
        .Y(n2681) );
  AOI2BB2X4 U2978 ( .B0(n2144), .B1(\U3/temp9t[6] ), .A0N(n2683), .A1N(n2674), 
        .Y(n2682) );
  AOI2BB2X4 U2979 ( .B0(n2144), .B1(\U3/temp9t[5] ), .A0N(n2690), .A1N(n2673), 
        .Y(n2683) );
  AOI2BB2X4 U2980 ( .B0(n2144), .B1(\U3/temp9t[4] ), .A0N(n2684), .A1N(n2672), 
        .Y(n2690) );
  AOI2BB2X4 U2981 ( .B0(n2144), .B1(\U3/temp9t[3] ), .A0N(n2671), .A1N(n2195), 
        .Y(n2684) );
  AOI2BB2X4 U2982 ( .B0(n2144), .B1(\U3/temp9t[2] ), .A0N(n2686), .A1N(n2194), 
        .Y(n2671) );
  OAI21X4 U2983 ( .A0(n2534), .A1(n2508), .B0(n2509), .Y(\U2/temp_x[11] ) );
  AOI2BB2X2 U2984 ( .B0(n2513), .B1(n738), .A0N(n738), .A1N(n2530), .Y(n2508)
         );
  AND3X4 U2985 ( .A(n2459), .B(n2460), .C(n2461), .Y(n2525) );
  NOR2BX4 U2986 ( .AN(n2432), .B(n2433), .Y(n2523) );
  AND3X4 U2987 ( .A(n2422), .B(n2421), .C(n2420), .Y(n2524) );
  AND3X4 U2988 ( .A(n2390), .B(n2391), .C(n2392), .Y(n1698) );
  AND2X4 U2989 ( .A(n2356), .B(n2357), .Y(n1700) );
  NOR2X4 U2990 ( .A(n751), .B(n725), .Y(n1709) );
  INVX8 U2991 ( .A(n1671), .Y(n732) );
  INVX8 U2992 ( .A(n2546), .Y(n731) );
  CLKINVX3 U2993 ( .A(n2516), .Y(n2519) );
  NAND2X1 U2994 ( .A(n966), .B(n1463), .Y(n2474) );
  NAND2X4 U2995 ( .A(n963), .B(n966), .Y(n2473) );
  NAND2X4 U2996 ( .A(n963), .B(n1463), .Y(n2472) );
  INVX8 U2997 ( .A(n2469), .Y(n963) );
  NAND2X4 U2998 ( .A(n2468), .B(n2467), .Y(n2469) );
  OAI21X4 U2999 ( .A0(n968), .A1(n1471), .B0(n2463), .Y(n2462) );
  AND3X4 U3000 ( .A(n2319), .B(n2318), .C(n2320), .Y(n1476) );
  OAI2BB1X4 U3001 ( .A0N(n966), .A1N(n1482), .B0(n2288), .Y(n1479) );
  NOR3X4 U3002 ( .A(n2285), .B(n2284), .C(n2283), .Y(n1482) );
  AND3X4 U3003 ( .A(n2347), .B(n2349), .C(n2348), .Y(n2535) );
  AND3X4 U3004 ( .A(n2205), .B(n2204), .C(n2203), .Y(n1870) );
  XOR2X4 U3005 ( .A(n1895), .B(n1896), .Y(n2544) );
  AND3X4 U3006 ( .A(n2181), .B(n2182), .C(n2183), .Y(n1875) );
  AOI2BB2X4 U3007 ( .B0(n1934), .B1(n2527), .A0N(n1934), .A1N(n2527), .Y(n1871) );
  XOR2X2 U3008 ( .A(n661), .B(n1912), .Y(n1934) );
  XNOR2X2 U3009 ( .A(n2550), .B(n660), .Y(n1891) );
  BUFX12 U3010 ( .A(n1859), .Y(n2547) );
  INVX8 U3011 ( .A(n2330), .Y(n1904) );
  INVX8 U3012 ( .A(n2238), .Y(n1906) );
  OAI222X4 U3013 ( .A0(n2527), .A1(n661), .B0(n2527), .B1(n1912), .C0(n661), 
        .C1(n1912), .Y(n1911) );
  OAI222X4 U3014 ( .A0(n1890), .A1(n2571), .B0(n1890), .B1(n2164), .C0(n2571), 
        .C1(n2164), .Y(n1894) );
  XOR2X4 U3015 ( .A(n1921), .B(n1922), .Y(n1909) );
  AOI21X4 U3016 ( .A0(n2578), .A1(n2590), .B0(n2577), .Y(n2165) );
  CLKINVX3 U3017 ( .A(n2184), .Y(n2577) );
  AOI222X4 U3018 ( .A0(n837), .A1(n1950), .B0(n837), .B1(n1947), .C0(n1947), 
        .C1(n1950), .Y(n1942) );
  AOI21X4 U3019 ( .A0(\U5/temp5t[0] ), .A1(\U5/U5/temp[0] ), .B0(n1400), .Y(
        n1389) );
  INVX8 U3020 ( .A(n2413), .Y(n1969) );
  BUFX12 U3021 ( .A(n1962), .Y(n2538) );
  AND3X4 U3022 ( .A(n2189), .B(n2188), .C(n2187), .Y(n1977) );
  INVX8 U3023 ( .A(n1987), .Y(n639) );
  OAI2BB2X4 U3024 ( .B0(n2032), .B1(n2583), .A0N(n2032), .A1N(n2583), .Y(n1987) );
  XNOR2X2 U3025 ( .A(n2587), .B(n2017), .Y(n2032) );
  INVX8 U3026 ( .A(n2554), .Y(n646) );
  OAI2BB1X4 U3027 ( .A0N(n2325), .A1N(n2324), .B0(n2326), .Y(n2011) );
  OR2X4 U3028 ( .A(n2269), .B(n2270), .Y(n2000) );
  OAI222X4 U3029 ( .A0(n1989), .A1(n1993), .B0(n1989), .B1(n1992), .C0(n1993), 
        .C1(n1992), .Y(n1998) );
  XOR2X4 U3030 ( .A(n2018), .B(n1914), .Y(n2014) );
  XNOR2X4 U3031 ( .A(n2184), .B(n2590), .Y(n1916) );
  XNOR2X4 U3032 ( .A(n835), .B(n1923), .Y(n1918) );
  NAND2X2 U3033 ( .A(n1930), .B(n1926), .Y(n2231) );
  XOR2X4 U3034 ( .A(n2035), .B(n1819), .Y(n1938) );
  CLKINVX3 U3035 ( .A(n1846), .Y(n2600) );
  NOR2X4 U3036 ( .A(n800), .B(n851), .Y(n1285) );
  INVX8 U3037 ( .A(n1432), .Y(n985) );
  XOR2X4 U3038 ( .A(n2506), .B(n2131), .Y(\U2/temp_y[11] ) );
  OAI21X4 U3039 ( .A0(n739), .A1(n726), .B0(n2507), .Y(n2506) );
  INVX8 U3040 ( .A(n1668), .Y(n726) );
  OAI21X4 U3041 ( .A0(n2545), .A1(n2129), .B0(n2504), .Y(n1668) );
  OAI22X4 U3042 ( .A0(n1637), .A1(n2484), .B0(n2530), .B1(n730), .Y(n1635) );
  OAI222X4 U3043 ( .A0(n2546), .A1(n739), .B0(n2546), .B1(n1640), .C0(n739), 
        .C1(n1640), .Y(n1637) );
  AOI2BB2X4 U3044 ( .B0(n1818), .B1(n1747), .A0N(n1818), .A1N(n1747), .Y(n1672) );
  XOR2X2 U3045 ( .A(n761), .B(n1771), .Y(n1818) );
  AND3X4 U3046 ( .A(n2441), .B(n2440), .C(n2442), .Y(n1653) );
  XNOR2X2 U3047 ( .A(n2434), .B(n1759), .Y(n1758) );
  XOR2X4 U3048 ( .A(n1760), .B(n1715), .Y(n1641) );
  XOR2X2 U3049 ( .A(n1716), .B(n740), .Y(n1760) );
  XOR2X4 U3050 ( .A(n1749), .B(n2400), .Y(n2401) );
  XOR2X2 U3051 ( .A(n2585), .B(n1751), .Y(n1749) );
  AND3X4 U3052 ( .A(n2384), .B(n2385), .C(n2386), .Y(n1751) );
  AND3X4 U3053 ( .A(n2362), .B(n2363), .C(n2364), .Y(n1725) );
  OAI222X4 U3054 ( .A0(n1732), .A1(n762), .B0(n1732), .B1(n2147), .C0(n762), 
        .C1(n2147), .Y(n1770) );
  OAI21X4 U3055 ( .A0(n1771), .A1(n761), .B0(n2218), .Y(n1733) );
  AND3X4 U3056 ( .A(n2173), .B(n2174), .C(n2175), .Y(n1683) );
  INVX8 U3057 ( .A(n1761), .Y(n740) );
  BUFX12 U3058 ( .A(n2427), .Y(n1750) );
  XOR2X4 U3059 ( .A(n1781), .B(n2135), .Y(n2309) );
  AND3X4 U3060 ( .A(n2397), .B(n2398), .C(n2399), .Y(n1757) );
  XOR2X4 U3061 ( .A(n1837), .B(n1823), .Y(n2219) );
  AND3X4 U3062 ( .A(n2299), .B(n2300), .C(n2301), .Y(n1745) );
  AOI222X4 U3063 ( .A0(n1735), .A1(n1684), .B0(n1735), .B1(n2146), .C0(n1684), 
        .C1(n2146), .Y(n1738) );
  XNOR2X4 U3064 ( .A(n1768), .B(n1769), .Y(n2157) );
  INVX8 U3065 ( .A(n2294), .Y(n1778) );
  INVX8 U3066 ( .A(n2336), .Y(n1772) );
  AOI21X4 U3067 ( .A0(n2586), .A1(n1834), .B0(n2286), .Y(n1805) );
  XNOR2X2 U3068 ( .A(n2581), .B(n2582), .Y(n2162) );
  INVX8 U3069 ( .A(n2126), .Y(n2563) );
  XNOR2X4 U3070 ( .A(n830), .B(n1765), .Y(n1788) );
  INVX8 U3071 ( .A(n1790), .Y(n772) );
  XOR2X4 U3072 ( .A(n1813), .B(n1812), .Y(n1790) );
  INVX8 U3073 ( .A(n2297), .Y(n2548) );
  XNOR2X2 U3074 ( .A(n1815), .B(n2143), .Y(n2290) );
  XOR2X2 U3075 ( .A(n1842), .B(n1822), .Y(n1803) );
  INVX8 U3076 ( .A(n2206), .Y(n2586) );
  XNOR2X4 U3077 ( .A(n1802), .B(n1801), .Y(n2159) );
  INVX8 U3078 ( .A(n2373), .Y(n1813) );
  NAND3BX4 U3079 ( .AN(n2372), .B(n2160), .C(n2371), .Y(n2373) );
  INVX8 U3080 ( .A(n2251), .Y(n1815) );
  OAI2BB2X4 U3081 ( .B0(n1040), .B1(temp1t[4]), .A0N(n1822), .A1N(n2250), .Y(
        n2251) );
  AND3X4 U3082 ( .A(n2167), .B(n2168), .C(n2169), .Y(n1822) );
  AND3X4 U3083 ( .A(n2196), .B(n2197), .C(n2198), .Y(n1841) );
  XOR2X1 U3084 ( .A(n2829), .B(n2737), .Y(n2714) );
  XOR2X1 U3085 ( .A(n2762), .B(n2761), .Y(\U3/Ytt[2] ) );
  XOR2X1 U3086 ( .A(n2760), .B(n2759), .Y(n2761) );
  AND2X2 U3087 ( .A(\intadd_25/SUM[8] ), .B(n2302), .Y(\intadd_51/B[0] ) );
  XOR2X1 U3088 ( .A(n1174), .B(n1175), .Y(temp5[8]) );
  AOI222X4 U3089 ( .A0(x3[6]), .A1(n618), .B0(x3[6]), .B1(n607), .C0(n618), 
        .C1(n607), .Y(n1176) );
  XOR2X1 U3090 ( .A(n1142), .B(n1143), .Y(temp7[8]) );
  AOI222X4 U3091 ( .A0(x1[6]), .A1(n628), .B0(x1[6]), .B1(n579), .C0(n628), 
        .C1(n579), .Y(n1144) );
  OAI2BB1X4 U3092 ( .A0N(n2828), .A1N(n2827), .B0(n2826), .Y(n2838) );
  AND2X2 U3093 ( .A(n2806), .B(\intadd_28/n1 ), .Y(n2803) );
  AND2X2 U3094 ( .A(\intadd_28/n1 ), .B(n2796), .Y(n2797) );
  OAI2BB1X4 U3095 ( .A0N(n2747), .A1N(n2754), .B0(n2746), .Y(n2798) );
  AND2X2 U3096 ( .A(n2736), .B(n2829), .Y(n2738) );
  AND2X2 U3097 ( .A(n2660), .B(n2658), .Y(n2659) );
  CLKINVX3 U3098 ( .A(n2756), .Y(n2745) );
  AND2X2 U3099 ( .A(\intadd_28/n1 ), .B(n2836), .Y(n2726) );
  INVX4 U3100 ( .A(n2702), .Y(n2732) );
  OAI2BB1X4 U3101 ( .A0N(n2701), .A1N(n2700), .B0(n2699), .Y(\intadd_28/n1 )
         );
  AND2X2 U3102 ( .A(n2836), .B(n2749), .Y(n2665) );
  AND2X2 U3103 ( .A(n2647), .B(n2730), .Y(n2648) );
  AND2X2 U3104 ( .A(n2730), .B(n2708), .Y(n2643) );
  XOR2X1 U3105 ( .A(n2641), .B(n2640), .Y(n2661) );
  XOR2X1 U3106 ( .A(\U3/temp12[12] ), .B(\U3/temp10t[2] ), .Y(n2640) );
  INVX8 U3107 ( .A(n2836), .Y(n2727) );
  AND2X2 U3108 ( .A(\U3/temp12[0] ), .B(n2607), .Y(n2639) );
  XOR2X1 U3109 ( .A(n2291), .B(n2842), .Y(n2818) );
  CLKINVX3 U3110 ( .A(n1210), .Y(n578) );
  AND2X2 U3111 ( .A(n1302), .B(n1323), .Y(n2448) );
  OAI222X4 U3112 ( .A0(n1313), .A1(n1302), .B0(n1313), .B1(n1006), .C0(n1302), 
        .C1(n1006), .Y(n1310) );
  AOI222X4 U3113 ( .A0(n1003), .A1(n1001), .B0(n1003), .B1(n1319), .C0(n1001), 
        .C1(n1319), .Y(n1315) );
  OAI222X4 U3114 ( .A0(n1306), .A1(n1322), .B0(n1306), .B1(n1005), .C0(n1322), 
        .C1(n1005), .Y(n1318) );
  AOI222X4 U3115 ( .A0(n1325), .A1(n2140), .B0(n1325), .B1(n1326), .C0(n2140), 
        .C1(n1326), .Y(n1321) );
  AOI222X4 U3116 ( .A0(n1008), .A1(n1072), .B0(n1008), .B1(n1337), .C0(n1072), 
        .C1(n1337), .Y(n1325) );
  XNOR2X2 U3117 ( .A(n1344), .B(n1351), .Y(n1327) );
  AOI222X4 U3118 ( .A0(\U5/U6/temp[11] ), .A1(n1335), .B0(\U5/U6/temp[11] ), 
        .B1(n1054), .C0(n1335), .C1(n1054), .Y(n1332) );
  AOI222X4 U3119 ( .A0(\U5/U6/temp[4] ), .A1(n1010), .B0(\U5/U6/temp[4] ), 
        .B1(n1344), .C0(n1010), .C1(n1344), .Y(n1335) );
  AOI222X4 U3120 ( .A0(\U5/U6/temp[6] ), .A1(n1349), .B0(\U5/U6/temp[6] ), 
        .B1(n1052), .C0(n1349), .C1(n1052), .Y(n1344) );
  AOI222X4 U3121 ( .A0(\U5/U6/temp[2] ), .A1(n1054), .B0(\U5/U6/temp[2] ), 
        .B1(n1341), .C0(n1054), .C1(n1341), .Y(n1349) );
  AOI222X4 U3122 ( .A0(\U5/U6/temp[4] ), .A1(n1328), .B0(\U5/U6/temp[4] ), 
        .B1(n1092), .C0(n1328), .C1(n1092), .Y(n1341) );
  AOI222X4 U3123 ( .A0(\U5/U6/temp[0] ), .A1(n1052), .B0(\U5/U6/temp[0] ), 
        .B1(n1339), .C0(n1052), .C1(n1339), .Y(n1328) );
  AOI222X4 U3124 ( .A0(\U5/U6/temp[2] ), .A1(n1333), .B0(\U5/U6/temp[2] ), 
        .B1(n1074), .C0(n1333), .C1(n1074), .Y(n1339) );
  AOI222X4 U3125 ( .A0(\U5/temp7t[1] ), .A1(n1092), .B0(\U5/temp7t[1] ), .B1(
        n1346), .C0(n1092), .C1(n1346), .Y(n1333) );
  XOR2X1 U3126 ( .A(n1292), .B(\intadd_42/n1 ), .Y(\U5/temp7[10] ) );
  MXI2X2 U3127 ( .A(n692), .B(\intadd_39/n1 ), .S0(n1284), .Y(\intadd_33/A[6] ) );
  OAI2BB2X2 U3128 ( .B0(\intadd_45/A[8] ), .B1(\intadd_39/B[8] ), .A0N(
        \intadd_39/B[8] ), .A1N(\intadd_45/A[8] ), .Y(n1284) );
  INVX8 U3129 ( .A(n1515), .Y(n691) );
  INVX8 U3130 ( .A(n1513), .Y(n690) );
  OAI222X4 U3131 ( .A0(\intadd_45/A[8] ), .A1(\intadd_39/B[8] ), .B0(
        \intadd_45/A[8] ), .B1(n694), .C0(\intadd_39/B[8] ), .C1(n694), .Y(
        n1513) );
  CLKINVX3 U3132 ( .A(n2057), .Y(n777) );
  OAI222X4 U3133 ( .A0(n692), .A1(\intadd_39/B[8] ), .B0(n692), .B1(n776), 
        .C0(\intadd_39/B[8] ), .C1(n776), .Y(n1515) );
  OAI21X4 U3134 ( .A0(n1296), .A1(n778), .B0(n1297), .Y(\intadd_45/A[8] ) );
  XOR2X2 U3135 ( .A(n1269), .B(n1270), .Y(\intadd_39/B[6] ) );
  AOI2BB2X2 U3136 ( .B0(n1245), .B1(n1246), .A0N(n1246), .A1N(n1245), .Y(n2055) );
  AOI2BB2X2 U3137 ( .B0(n1278), .B1(n1270), .A0N(n1270), .A1N(n1278), .Y(n2056) );
  OAI21X4 U3138 ( .A0(n1294), .A1(n1268), .B0(n1295), .Y(\intadd_39/B[8] ) );
  AOI222X4 U3139 ( .A0(n1056), .A1(n1013), .B0(n1056), .B1(n1269), .C0(n1013), 
        .C1(n1269), .Y(n1268) );
  OAI222X4 U3140 ( .A0(n1094), .A1(n1060), .B0(n1094), .B1(n1272), .C0(n1060), 
        .C1(n1272), .Y(n1271) );
  OAI222X4 U3141 ( .A0(n1274), .A1(\U5/temp1[4] ), .B0(n1274), .B1(
        \U5/temp2[4] ), .C0(\U5/temp1[4] ), .C1(\U5/temp2[4] ), .Y(n1272) );
  OAI222X4 U3142 ( .A0(n1111), .A1(n1100), .B0(n1111), .B1(n1275), .C0(n1100), 
        .C1(n1275), .Y(n1274) );
  OAI222X4 U3143 ( .A0(n720), .A1(\U5/temp1[2] ), .B0(n720), .B1(\U5/temp2[2] ), .C0(\U5/temp1[2] ), .C1(\U5/temp2[2] ), .Y(n1275) );
  OAI222X4 U3144 ( .A0(n1056), .A1(\U5/temp2[7] ), .B0(n1056), .B1(n1278), 
        .C0(\U5/temp2[7] ), .C1(n1278), .Y(n1243) );
  OAI222X4 U3145 ( .A0(n1097), .A1(\U5/temp1[6] ), .B0(n1097), .B1(n1245), 
        .C0(\U5/temp1[6] ), .C1(n1245), .Y(n1278) );
  OAI222X4 U3146 ( .A0(n1094), .A1(\U5/temp2[5] ), .B0(n1094), .B1(n1279), 
        .C0(\U5/temp2[5] ), .C1(n1279), .Y(n1245) );
  OAI222X4 U3147 ( .A0(n1096), .A1(\U5/temp1[4] ), .B0(n1096), .B1(n1247), 
        .C0(\U5/temp1[4] ), .C1(n1247), .Y(n1279) );
  OAI222X4 U3148 ( .A0(n1111), .A1(\U5/temp2[3] ), .B0(n1111), .B1(n1280), 
        .C0(\U5/temp2[3] ), .C1(n1280), .Y(n1247) );
  OAI222X4 U3149 ( .A0(n1125), .A1(\U5/temp1[2] ), .B0(n1125), .B1(n785), .C0(
        \U5/temp1[2] ), .C1(n785), .Y(n1280) );
  MXI2X2 U3150 ( .A(n992), .B(n1354), .S0(n2453), .Y(\U5/Xt[8] ) );
  AOI2BB2X2 U3151 ( .B0(n2536), .B1(n1957), .A0N(n2536), .A1N(n1957), .Y(n2501) );
  AOI2BB2X2 U3152 ( .B0(n2536), .B1(n640), .A0N(n2536), .A1N(n640), .Y(n2500)
         );
  AOI2BB2X4 U3153 ( .B0(n2415), .B1(n2416), .A0N(n2816), .A1N(n2839), .Y(n2822) );
  INVX8 U3154 ( .A(n2409), .Y(n2816) );
  AOI21X4 U3155 ( .A0(n2406), .A1(n2785), .B0(n2408), .Y(n2409) );
  AOI2BB2X4 U3156 ( .B0(n2395), .B1(n2786), .A0N(n2789), .A1N(n2396), .Y(n2785) );
  OAI2BB1X4 U3157 ( .A0N(n2393), .A1N(n2777), .B0(n2394), .Y(n2792) );
  NOR2BX4 U3158 ( .AN(n2381), .B(n2382), .Y(n2777) );
  XOR2X1 U3159 ( .A(n2210), .B(n2773), .Y(n2774) );
  OAI2BB1X4 U3160 ( .A0N(n2768), .A1N(n2771), .B0(n2767), .Y(n2787) );
  AOI2BB2X4 U3161 ( .B0(n2842), .B1(n2233), .A0N(n2295), .A1N(n2246), .Y(n2771) );
  AND2X2 U3162 ( .A(n2840), .B(n2842), .Y(n2475) );
  AND2X2 U3163 ( .A(n2770), .B(n2813), .Y(n2296) );
  AND2X2 U3164 ( .A(n2202), .B(n2210), .Y(n2224) );
  CLKINVX3 U3165 ( .A(n2688), .Y(n2773) );
  AND2X2 U3166 ( .A(n2689), .B(n2670), .Y(n2687) );
  XOR2X1 U3167 ( .A(\U3/temp9t[2] ), .B(n2144), .Y(n2685) );
  AOI2BB2X4 U3168 ( .B0(\U3/temp12[1] ), .B1(n2144), .A0N(n2696), .A1N(n2695), 
        .Y(n2716) );
  XOR2X1 U3169 ( .A(n2146), .B(n1735), .Y(n1734) );
  AND3X4 U3170 ( .A(n2472), .B(n2473), .C(n2474), .Y(n1461) );
  OAI222X4 U3171 ( .A0(n1474), .A1(n1463), .B0(n1474), .B1(n970), .C0(n1463), 
        .C1(n970), .Y(n1471) );
  OAI2BB1X2 U3172 ( .A0N(n1493), .A1N(\U4/U5/temp[6] ), .B0(n2268), .Y(n2266)
         );
  AND2X2 U3173 ( .A(n973), .B(n1487), .Y(n2283) );
  XNOR2X2 U3174 ( .A(n1496), .B(n2185), .Y(n1484) );
  XNOR2X2 U3175 ( .A(n1505), .B(n1512), .Y(n1488) );
  AOI21X4 U3176 ( .A0(\U4/temp5t[0] ), .A1(\U4/U5/temp[0] ), .B0(n1509), .Y(
        n1498) );
  XNOR2X4 U3177 ( .A(n1493), .B(n1504), .Y(n1467) );
  INVX8 U3178 ( .A(n1463), .Y(n968) );
  AOI222X4 U3179 ( .A0(\U4/U5/temp[11] ), .A1(n1496), .B0(\U4/U5/temp[11] ), 
        .B1(n1045), .C0(n1496), .C1(n1045), .Y(n1493) );
  AOI222X4 U3180 ( .A0(\U4/U5/temp[4] ), .A1(n974), .B0(\U4/U5/temp[4] ), .B1(
        n1505), .C0(n974), .C1(n1505), .Y(n1496) );
  AOI222X4 U3181 ( .A0(\U4/U5/temp[6] ), .A1(n1510), .B0(\U4/U5/temp[6] ), 
        .B1(n1043), .C0(n1510), .C1(n1043), .Y(n1505) );
  AOI222X4 U3182 ( .A0(\U4/U5/temp[2] ), .A1(n1045), .B0(\U4/U5/temp[2] ), 
        .B1(n1502), .C0(n1045), .C1(n1502), .Y(n1510) );
  AOI222X4 U3183 ( .A0(\U4/U5/temp[4] ), .A1(n1489), .B0(\U4/U5/temp[4] ), 
        .B1(n1086), .C0(n1489), .C1(n1086), .Y(n1502) );
  AOI222X4 U3184 ( .A0(\U4/U5/temp[0] ), .A1(n1043), .B0(\U4/U5/temp[0] ), 
        .B1(n1500), .C0(n1043), .C1(n1500), .Y(n1489) );
  AOI222X4 U3185 ( .A0(\U4/U5/temp[2] ), .A1(n1494), .B0(\U4/U5/temp[2] ), 
        .B1(n1066), .C0(n1494), .C1(n1066), .Y(n1500) );
  AOI222X4 U3186 ( .A0(\U4/temp5t[1] ), .A1(n1086), .B0(\U4/temp5t[1] ), .B1(
        n1507), .C0(n1086), .C1(n1507), .Y(n1494) );
  CLKINVX3 U3187 ( .A(n1867), .Y(n659) );
  AND3X4 U3188 ( .A(n2260), .B(n2261), .C(n2262), .Y(n1868) );
  XOR2X2 U3189 ( .A(n671), .B(n1897), .Y(n1895) );
  AOI222X4 U3190 ( .A0(n1867), .A1(n1880), .B0(n1867), .B1(n1881), .C0(n1880), 
        .C1(n1881), .Y(n1878) );
  NOR2X4 U3191 ( .A(n1871), .B(n1933), .Y(n1881) );
  XOR2X1 U3192 ( .A(n1893), .B(n1894), .Y(n1892) );
  AOI2BB2X2 U3193 ( .B0(n1898), .B1(n2540), .A0N(n1898), .A1N(n2540), .Y(n1865) );
  XOR2X2 U3194 ( .A(n2527), .B(n1901), .Y(n1898) );
  INVX8 U3195 ( .A(n2549), .Y(n654) );
  OAI2BB1X4 U3196 ( .A0N(n668), .A1N(n1904), .B0(n1903), .Y(n2374) );
  AOI222X4 U3197 ( .A0(n1919), .A1(n1920), .B0(n1919), .B1(n1921), .C0(n1920), 
        .C1(n1921), .Y(n1903) );
  AND2X4 U3198 ( .A(n2275), .B(n2274), .Y(n1908) );
  INVX8 U3199 ( .A(n1910), .Y(n671) );
  AOI222X4 U3200 ( .A0(n670), .A1(n2527), .B0(n670), .B1(n1901), .C0(n1901), 
        .C1(n2527), .Y(n1897) );
  AND3X4 U3201 ( .A(n2180), .B(n2179), .C(n2178), .Y(n1901) );
  OAI222X4 U3202 ( .A0(n1887), .A1(n1886), .B0(n1886), .B1(n2550), .C0(n1887), 
        .C1(n2550), .Y(n1912) );
  OAI222X4 U3203 ( .A0(n1943), .A1(n677), .B0(n1943), .B1(n1894), .C0(n677), 
        .C1(n1894), .Y(n1887) );
  XOR2X2 U3204 ( .A(n1929), .B(n1935), .Y(n1900) );
  AND3X4 U3205 ( .A(n2241), .B(n2243), .C(n2242), .Y(n1921) );
  NAND2X2 U3206 ( .A(n1917), .B(n835), .Y(n2241) );
  NOR2X4 U3207 ( .A(n2165), .B(n2166), .Y(n1917) );
  NOR2X4 U3208 ( .A(n2578), .B(n2590), .Y(n2166) );
  AOI222X4 U3209 ( .A0(n1926), .A1(n836), .B0(n1926), .B1(n1913), .C0(n1913), 
        .C1(n836), .Y(n1915) );
  AOI222X4 U3210 ( .A0(n1927), .A1(n1928), .B0(n1927), .B1(n1929), .C0(n1928), 
        .C1(n1929), .Y(n1913) );
  AOI222X4 U3211 ( .A0(n832), .A1(n1936), .B0(n832), .B1(n1937), .C0(n1937), 
        .C1(n1936), .Y(n1929) );
  AOI222X4 U3212 ( .A0(n1940), .A1(n2125), .B0(n1940), .B1(n2589), .C0(n2125), 
        .C1(n2589), .Y(n1937) );
  AOI222X4 U3213 ( .A0(n1953), .A1(n1954), .B0(n1953), .B1(n2564), .C0(n1954), 
        .C1(n2564), .Y(n1945) );
  AND3X4 U3214 ( .A(n2490), .B(n2491), .C(n2492), .Y(n1959) );
  AND2X2 U3215 ( .A(n1354), .B(n1375), .Y(n2428) );
  OAI222X4 U3216 ( .A0(n1365), .A1(n1354), .B0(n1365), .B1(n994), .C0(n1354), 
        .C1(n994), .Y(n1362) );
  OAI222X4 U3217 ( .A0(n992), .A1(n1368), .B0(n992), .B1(n988), .C0(n1368), 
        .C1(n988), .Y(n1365) );
  AOI222X4 U3218 ( .A0(\U5/U5/temp[6] ), .A1(n1021), .B0(\U5/U5/temp[6] ), 
        .B1(n1384), .C0(n1021), .C1(n1384), .Y(n1382) );
  AOI222X4 U3219 ( .A0(n1377), .A1(n997), .B0(n1377), .B1(n1378), .C0(n997), 
        .C1(n1378), .Y(n1373) );
  AOI222X4 U3220 ( .A0(n996), .A1(n1077), .B0(n996), .B1(n1389), .C0(n1077), 
        .C1(n1389), .Y(n1377) );
  INVX8 U3221 ( .A(n1354), .Y(n992) );
  AOI222X4 U3222 ( .A0(\U5/U5/temp[11] ), .A1(n1387), .B0(\U5/U5/temp[11] ), 
        .B1(n1051), .C0(n1387), .C1(n1051), .Y(n1384) );
  AOI222X4 U3223 ( .A0(\U5/U5/temp[4] ), .A1(n998), .B0(\U5/U5/temp[4] ), .B1(
        n1396), .C0(n998), .C1(n1396), .Y(n1387) );
  AOI222X4 U3224 ( .A0(\U5/U5/temp[6] ), .A1(n1401), .B0(\U5/U5/temp[6] ), 
        .B1(n1049), .C0(n1401), .C1(n1049), .Y(n1396) );
  AOI222X4 U3225 ( .A0(\U5/U5/temp[2] ), .A1(n1051), .B0(\U5/U5/temp[2] ), 
        .B1(n1393), .C0(n1051), .C1(n1393), .Y(n1401) );
  AOI222X4 U3226 ( .A0(\U5/U5/temp[4] ), .A1(n1380), .B0(\U5/U5/temp[4] ), 
        .B1(n1090), .C0(n1380), .C1(n1090), .Y(n1393) );
  AOI222X4 U3227 ( .A0(\U5/U5/temp[0] ), .A1(n1049), .B0(\U5/U5/temp[0] ), 
        .B1(n1391), .C0(n1049), .C1(n1391), .Y(n1380) );
  AOI222X4 U3228 ( .A0(\U5/U5/temp[2] ), .A1(n1385), .B0(\U5/U5/temp[2] ), 
        .B1(n1071), .C0(n1385), .C1(n1071), .Y(n1391) );
  AOI222X4 U3229 ( .A0(\U5/temp5t[1] ), .A1(n1090), .B0(\U5/temp5t[1] ), .B1(
        n1398), .C0(n1090), .C1(n1398), .Y(n1385) );
  AND3X4 U3230 ( .A(n2464), .B(n2465), .C(n2466), .Y(n1961) );
  AND3X4 U3231 ( .A(n2438), .B(n2437), .C(n2439), .Y(n1965) );
  AND3X4 U3232 ( .A(n2429), .B(n2430), .C(n2431), .Y(n1968) );
  XOR2X4 U3233 ( .A(n2001), .B(n2379), .Y(n2380) );
  XOR2X2 U3234 ( .A(n2127), .B(n2004), .Y(n2001) );
  AND3X4 U3235 ( .A(n2387), .B(n2388), .C(n2389), .Y(n1973) );
  OAI222X4 U3236 ( .A0(n646), .A1(n638), .B0(n646), .B1(n1983), .C0(n638), 
        .C1(n1983), .Y(n1981) );
  CLKINVX3 U3237 ( .A(n2532), .Y(n2583) );
  AOI2BB2X4 U3238 ( .B0(n2005), .B1(n666), .A0N(n2005), .A1N(n666), .Y(n2579)
         );
  AOI31X4 U3239 ( .A0(n664), .A1(n2333), .A2(n2004), .B0(n2002), .Y(n1957) );
  OAI222X4 U3240 ( .A0(n1920), .A1(n672), .B0(n1920), .B1(n665), .C0(n672), 
        .C1(n665), .Y(n2002) );
  OAI2BB1X4 U3241 ( .A0N(n666), .A1N(n2367), .B0(n2365), .Y(n2004) );
  OAI222X4 U3242 ( .A0(n2014), .A1(n1995), .B0(n2014), .B1(n662), .C0(n662), 
        .C1(n1995), .Y(n2007) );
  OAI222X4 U3243 ( .A0(n663), .A1(n2016), .B0(n2017), .B1(n2016), .C0(n2017), 
        .C1(n663), .Y(n1995) );
  OAI222X4 U3244 ( .A0(n2015), .A1(n1990), .B0(n2015), .B1(n674), .C0(n1990), 
        .C1(n674), .Y(n2017) );
  XOR2X2 U3245 ( .A(n1935), .B(n2026), .Y(n2006) );
  INVX8 U3246 ( .A(n2161), .Y(n666) );
  XOR2X4 U3247 ( .A(n2019), .B(n1916), .Y(n2161) );
  INVX8 U3248 ( .A(n2020), .Y(n665) );
  AOI222X4 U3249 ( .A0(n1923), .A1(n2021), .B0(n1923), .B1(n1931), .C0(n2021), 
        .C1(n1931), .Y(n2020) );
  XOR2X4 U3250 ( .A(n2022), .B(n1796), .Y(n1931) );
  AOI222X4 U3251 ( .A0(temp2t[8]), .A1(temp3t[8]), .B0(temp2t[8]), .B1(n2024), 
        .C0(temp3t[8]), .C1(n2024), .Y(n2022) );
  AOI222X4 U3252 ( .A0(n2590), .A1(n2184), .B0(n2590), .B1(n2019), .C0(n2184), 
        .C1(n2019), .Y(n2021) );
  AND3X4 U3253 ( .A(n2229), .B(n2230), .C(n2231), .Y(n2019) );
  XOR2X4 U3254 ( .A(n2025), .B(n1799), .Y(n1930) );
  XOR2X4 U3255 ( .A(n2027), .B(n1801), .Y(n1926) );
  AND3X4 U3256 ( .A(n2215), .B(n2216), .C(n2217), .Y(n2018) );
  XOR2X4 U3257 ( .A(n2030), .B(n1808), .Y(n1927) );
  AOI222X4 U3258 ( .A0(n1936), .A1(n2033), .B0(n1936), .B1(n1938), .C0(n2033), 
        .C1(n1938), .Y(n2026) );
  AOI222X4 U3259 ( .A0(n831), .A1(n2125), .B0(n831), .B1(n2040), .C0(n2125), 
        .C1(n2040), .Y(n2033) );
  AOI222X4 U3260 ( .A0(n1950), .A1(n2036), .B0(n1950), .B1(n1956), .C0(n2036), 
        .C1(n1956), .Y(n2040) );
  AOI222X4 U3261 ( .A0(n838), .A1(n1952), .B0(n838), .B1(n2037), .C0(n1952), 
        .C1(n2037), .Y(n2036) );
  CLKINVX3 U3262 ( .A(n1842), .Y(n2573) );
  CLKINVX3 U3263 ( .A(n1940), .Y(n831) );
  INVX8 U3264 ( .A(n2591), .Y(n1936) );
  XOR2X2 U3265 ( .A(n2034), .B(n2143), .Y(n2591) );
  XOR2X4 U3266 ( .A(n673), .B(n1812), .Y(n2184) );
  OAI222X4 U3267 ( .A0(n2027), .A1(temp4t[7]), .B0(n2027), .B1(temp1t[7]), 
        .C0(temp4t[7]), .C1(temp1t[7]), .Y(n2028) );
  OAI222X4 U3268 ( .A0(n1033), .A1(n1042), .B0(n1033), .B1(n2029), .C0(n1042), 
        .C1(n2029), .Y(n2027) );
  OAI222X4 U3269 ( .A0(n2034), .A1(temp1t[5]), .B0(n2034), .B1(temp4t[5]), 
        .C0(temp1t[5]), .C1(temp4t[5]), .Y(n2029) );
  OAI222X4 U3270 ( .A0(n1032), .A1(n1040), .B0(n1032), .B1(n2038), .C0(n1040), 
        .C1(n2038), .Y(n2034) );
  OAI222X4 U3271 ( .A0(n2046), .A1(temp1t[3]), .B0(n2046), .B1(temp4t[3]), 
        .C0(temp1t[3]), .C1(temp4t[3]), .Y(n2038) );
  OAI222X4 U3272 ( .A0(n1079), .A1(n1084), .B0(n1079), .B1(n2044), .C0(n1084), 
        .C1(n2044), .Y(n2046) );
  OAI222X4 U3273 ( .A0(temp1t[1]), .A1(temp4t[1]), .B0(temp1t[1]), .B1(n2567), 
        .C0(temp4t[1]), .C1(n2567), .Y(n2044) );
  AOI222X4 U3274 ( .A0(n2025), .A1(n1037), .B0(n2025), .B1(n1039), .C0(n1037), 
        .C1(n1039), .Y(n2024) );
  AOI222X4 U3275 ( .A0(temp2t[6]), .A1(temp3t[6]), .B0(temp2t[6]), .B1(n2030), 
        .C0(temp3t[6]), .C1(n2030), .Y(n2025) );
  AOI222X4 U3276 ( .A0(n2035), .A1(n1035), .B0(n2035), .B1(n1038), .C0(n1035), 
        .C1(n1038), .Y(n2030) );
  AOI222X4 U3277 ( .A0(temp2t[4]), .A1(temp3t[4]), .B0(temp2t[4]), .B1(n2039), 
        .C0(temp3t[4]), .C1(n2039), .Y(n2035) );
  AOI222X4 U3278 ( .A0(n2041), .A1(n1081), .B0(n2041), .B1(n1083), .C0(n1081), 
        .C1(n1083), .Y(n2039) );
  AOI222X4 U3279 ( .A0(temp2t[2]), .A1(temp3t[2]), .B0(temp2t[2]), .B1(n2045), 
        .C0(temp3t[2]), .C1(n2045), .Y(n2041) );
  AOI222X4 U3280 ( .A0(n1121), .A1(n1122), .B0(n1121), .B1(n2043), .C0(n1122), 
        .C1(n2043), .Y(n2045) );
  OAI222X4 U3281 ( .A0(n1422), .A1(n1411), .B0(n1422), .B1(n982), .C0(n1411), 
        .C1(n982), .Y(n1419) );
  AOI222X4 U3282 ( .A0(n979), .A1(n977), .B0(n979), .B1(n1428), .C0(n977), 
        .C1(n1428), .Y(n1424) );
  XOR2X2 U3283 ( .A(n1439), .B(n1440), .Y(n1412) );
  AOI222X4 U3284 ( .A0(\U4/U6/temp[6] ), .A1(n1020), .B0(\U4/U6/temp[6] ), 
        .B1(n1441), .C0(n1020), .C1(n1441), .Y(n1439) );
  AOI222X4 U3285 ( .A0(n2163), .A1(n985), .B0(n2163), .B1(n1435), .C0(n985), 
        .C1(n1435), .Y(n1430) );
  AND3X4 U3286 ( .A(n2352), .B(n2350), .C(n2351), .Y(n2163) );
  AND2X4 U3287 ( .A(n982), .B(n2186), .Y(n2543) );
  XOR2X1 U3288 ( .A(\U4/U6/temp[0] ), .B(\U4/temp7t[0] ), .Y(n2186) );
  XOR2X2 U3289 ( .A(n1458), .B(n1459), .Y(n1421) );
  INVX8 U3290 ( .A(n1411), .Y(n980) );
  AOI222X4 U3291 ( .A0(\U4/U6/temp[11] ), .A1(n1444), .B0(\U4/U6/temp[11] ), 
        .B1(n1048), .C0(n1444), .C1(n1048), .Y(n1441) );
  AOI222X4 U3292 ( .A0(\U4/U6/temp[4] ), .A1(n986), .B0(\U4/U6/temp[4] ), .B1(
        n1453), .C0(n986), .C1(n1453), .Y(n1444) );
  AOI222X4 U3293 ( .A0(\U4/U6/temp[6] ), .A1(n1458), .B0(\U4/U6/temp[6] ), 
        .B1(n1046), .C0(n1458), .C1(n1046), .Y(n1453) );
  AOI222X4 U3294 ( .A0(\U4/U6/temp[2] ), .A1(n1048), .B0(\U4/U6/temp[2] ), 
        .B1(n1450), .C0(n1048), .C1(n1450), .Y(n1458) );
  AOI222X4 U3295 ( .A0(\U4/U6/temp[4] ), .A1(n1437), .B0(\U4/U6/temp[4] ), 
        .B1(n1088), .C0(n1437), .C1(n1088), .Y(n1450) );
  AOI222X4 U3296 ( .A0(\U4/U6/temp[0] ), .A1(n1046), .B0(\U4/U6/temp[0] ), 
        .B1(n1448), .C0(n1046), .C1(n1448), .Y(n1437) );
  AOI222X4 U3297 ( .A0(\U4/U6/temp[2] ), .A1(n1442), .B0(\U4/U6/temp[2] ), 
        .B1(n1069), .C0(n1442), .C1(n1069), .Y(n1448) );
  AOI222X4 U3298 ( .A0(\U4/temp7t[1] ), .A1(n1088), .B0(\U4/temp7t[1] ), .B1(
        n1455), .C0(n1088), .C1(n1455), .Y(n1442) );
  AOI31X4 U3299 ( .A0(n2434), .A1(n1721), .A2(n1713), .B0(n1763), .Y(n1762) );
  AND3X4 U3300 ( .A(n2402), .B(n2403), .C(n2404), .Y(n1721) );
  OAI222X4 U3301 ( .A0(n1641), .A1(n1643), .B0(n1641), .B1(n1671), .C0(n1643), 
        .C1(n1671), .Y(n1640) );
  OAI222X4 U3302 ( .A0(n1644), .A1(n734), .B0(n1644), .B1(n1647), .C0(n734), 
        .C1(n1647), .Y(n1643) );
  OAI222X4 U3303 ( .A0(n1650), .A1(n2558), .B0(n1650), .B1(n1672), .C0(n2558), 
        .C1(n1672), .Y(n1647) );
  XOR2X2 U3304 ( .A(n1756), .B(n2537), .Y(n1648) );
  CLKINVX3 U3305 ( .A(n1741), .Y(n2435) );
  XOR2X4 U3306 ( .A(n1758), .B(n2126), .Y(n1644) );
  AOI222X4 U3307 ( .A0(n759), .A1(n2566), .B0(n759), .B1(n1680), .C0(n2566), 
        .C1(n1680), .Y(n1676) );
  AOI31X4 U3308 ( .A0(n1715), .A1(n740), .A2(n1716), .B0(n1717), .Y(n1714) );
  AOI222X4 U3309 ( .A0(n830), .A1(n1765), .B0(n830), .B1(n1795), .C0(n1765), 
        .C1(n1795), .Y(n1716) );
  AOI222X4 U3310 ( .A0(n2563), .A1(n2434), .B0(n2563), .B1(n1759), .C0(n2434), 
        .C1(n1759), .Y(n1761) );
  AOI222X4 U3311 ( .A0(n1757), .A1(n2537), .B0(n1757), .B1(n1750), .C0(n2537), 
        .C1(n1750), .Y(n1759) );
  AOI222X4 U3312 ( .A0(n1753), .A1(n1741), .B0(n1753), .B1(n1732), .C0(n1741), 
        .C1(n1732), .Y(n1755) );
  XOR2X4 U3313 ( .A(n1778), .B(n1769), .Y(n1741) );
  AOI222X4 U3314 ( .A0(n2553), .A1(n1747), .B0(n2553), .B1(n1748), .C0(n1747), 
        .C1(n1748), .Y(n1753) );
  NAND2X4 U3315 ( .A(n752), .B(n2566), .Y(n1730) );
  BUFX3 U3316 ( .A(n2569), .Y(n2584) );
  AOI222X4 U3317 ( .A0(n1785), .A1(n1786), .B0(n1785), .B1(n1787), .C0(n1786), 
        .C1(n1787), .Y(n1795) );
  AND3X4 U3318 ( .A(n2311), .B(n2312), .C(n2313), .Y(n1785) );
  AND3X4 U3319 ( .A(n2376), .B(n2377), .C(n2378), .Y(n1783) );
  AND3X4 U3320 ( .A(n2355), .B(n2354), .C(n2353), .Y(n1776) );
  CLKINVX3 U3321 ( .A(n1829), .Y(n2191) );
  XOR2X4 U3322 ( .A(n754), .B(n1788), .Y(n1715) );
  INVX8 U3323 ( .A(n1764), .Y(n830) );
  AOI222X4 U3324 ( .A0(n1764), .A1(n754), .B0(n1764), .B1(n1765), .C0(n754), 
        .C1(n1765), .Y(n1713) );
  OAI222X4 U3325 ( .A0(n1011), .A1(temp1t[9]), .B0(n1011), .B1(n771), .C0(
        temp1t[9]), .C1(n771), .Y(n1765) );
  AOI222X4 U3326 ( .A0(n770), .A1(n1787), .B0(n770), .B1(n1766), .C0(n1787), 
        .C1(n1766), .Y(n1789) );
  AOI222X4 U3327 ( .A0(n2528), .A1(n1781), .B0(n2528), .B1(n772), .C0(n1781), 
        .C1(n772), .Y(n1766) );
  AOI222X4 U3328 ( .A0(n773), .A1(n1780), .B0(n773), .B1(n1768), .C0(n1780), 
        .C1(n1768), .Y(n1781) );
  AND3X4 U3329 ( .A(n2263), .B(n2264), .C(n2265), .Y(n1768) );
  INVX8 U3330 ( .A(n2341), .Y(n1777) );
  AND3X4 U3331 ( .A(n2252), .B(n2253), .C(n2254), .Y(n1774) );
  AOI222X4 U3332 ( .A0(n2128), .A1(n1823), .B0(n2128), .B1(n768), .C0(n1823), 
        .C1(n768), .Y(n1793) );
  AOI22X2 U3333 ( .A0(temp1t[4]), .A1(temp4t[4]), .B0(n1040), .B1(n1032), .Y(
        n1842) );
  AOI222X4 U3334 ( .A0(n767), .A1(n2124), .B0(n767), .B1(n1824), .C0(n2124), 
        .C1(n1824), .Y(n1823) );
  AOI222X4 U3335 ( .A0(n2559), .A1(n1826), .B0(n2559), .B1(n1829), .C0(n1826), 
        .C1(n1829), .Y(n1830) );
  INVX8 U3336 ( .A(n2569), .Y(n1826) );
  INVX8 U3337 ( .A(n2370), .Y(n1780) );
  INVX8 U3338 ( .A(n2304), .Y(n1787) );
  XOR2X4 U3339 ( .A(n771), .B(n1798), .Y(n1786) );
  INVX8 U3340 ( .A(n1814), .Y(n771) );
  AOI222X4 U3341 ( .A0(temp4t[8]), .A1(n1813), .B0(temp4t[8]), .B1(n960), .C0(
        n1813), .C1(n960), .Y(n1814) );
  AND3X4 U3342 ( .A(n2279), .B(n2280), .C(n2281), .Y(n1807) );
  AOI222X4 U3343 ( .A0(temp4t[2]), .A1(n1847), .B0(temp4t[2]), .B1(n1079), 
        .C0(n1847), .C1(n1079), .Y(n1843) );
  AOI222X4 U3344 ( .A0(temp1t[1]), .A1(n1124), .B0(temp1t[1]), .B1(n787), .C0(
        n1124), .C1(n787), .Y(n1847) );
  INVX8 U3345 ( .A(n2551), .Y(n787) );
  NOR2X4 U3346 ( .A(n800), .B(n2541), .Y(n1282) );
  AOI222X4 U3347 ( .A0(temp3t[9]), .A1(n1012), .B0(temp3t[9]), .B1(n1797), 
        .C0(n1012), .C1(n1797), .Y(n1764) );
  AOI222X4 U3348 ( .A0(temp3t[8]), .A1(n1811), .B0(temp3t[8]), .B1(n961), .C0(
        n1811), .C1(n961), .Y(n1797) );
  AOI222X4 U3349 ( .A0(temp2t[7]), .A1(n1039), .B0(temp2t[7]), .B1(n2276), 
        .C0(n1039), .C1(n2276), .Y(n1811) );
  AND3X4 U3350 ( .A(n2255), .B(n2256), .C(n2257), .Y(n1816) );
  AND3X4 U3351 ( .A(n2207), .B(n2208), .C(n2209), .Y(n1820) );
  AOI222X4 U3352 ( .A0(temp2t[1]), .A1(n1122), .B0(temp2t[1]), .B1(n2542), 
        .C0(n1122), .C1(n2542), .Y(n1845) );
  XNOR3X2 U3353 ( .A(n2144), .B(\U3/temp11[1] ), .C(n2700), .Y(n2702) );
  INVX1 U3354 ( .A(\U3/temp10t[0] ), .Y(n2607) );
  XNOR3X2 U3355 ( .A(\U3/temp12[1] ), .B(n2606), .C(n2696), .Y(n2766) );
  AOI222X4 U3356 ( .A0(temp3t[9]), .A1(temp2t[9]), .B0(temp3t[9]), .B1(n2022), 
        .C0(temp2t[9]), .C1(n2022), .Y(n1920) );
  AOI222X4 U3357 ( .A0(temp4t[9]), .A1(temp1t[9]), .B0(temp4t[9]), .B1(n2023), 
        .C0(temp1t[9]), .C1(n2023), .Y(n1919) );
  AOI222X4 U3358 ( .A0(temp4t[8]), .A1(temp1t[8]), .B0(temp4t[8]), .B1(n673), 
        .C0(temp1t[8]), .C1(n673), .Y(n2023) );
  AOI21X1 U3359 ( .A0(n1871), .A1(n1933), .B0(n1881), .Y(n1932) );
  AOI2BB1X1 U3360 ( .A0N(\U1/result6[0] ), .A1N(\U1/temp_yyyt[0] ), .B0(
        \intadd_26/CI ), .Y(n2303) );
  AOI2BB1X1 U3361 ( .A0N(\U1/result5[0] ), .A1N(\U1/temp_xxxt[0] ), .B0(
        \intadd_25/CI ), .Y(n2302) );
  OAI21XL U3362 ( .A0(x4[8]), .A1(x3[8]), .B0(n1191), .Y(n1190) );
  INVX1 U3363 ( .A(n2759), .Y(n2740) );
  XNOR3X2 U3364 ( .A(n2709), .B(n2708), .C(n2707), .Y(n2737) );
  NAND2X1 U3365 ( .A(n2657), .B(n2656), .Y(n2658) );
  INVX1 U3366 ( .A(n2655), .Y(n2656) );
  XNOR3X2 U3367 ( .A(n2661), .B(n2734), .C(n2660), .Y(n2711) );
  XNOR3X2 U3368 ( .A(n2735), .B(n2734), .C(n2733), .Y(n2759) );
  XNOR3X2 U3369 ( .A(n2750), .B(n2730), .C(n2729), .Y(n2755) );
  NAND2X1 U3370 ( .A(n2702), .B(n2795), .Y(n2706) );
  OR2X2 U3371 ( .A(\intadd_28/n1 ), .B(n2752), .Y(n2747) );
  XNOR3X2 U3372 ( .A(n2794), .B(n2725), .C(n2724), .Y(n2752) );
  XNOR3X2 U3373 ( .A(n2750), .B(n2749), .C(n2748), .Y(n2796) );
  XNOR3X2 U3374 ( .A(n2795), .B(n2794), .C(n2793), .Y(n2809) );
  INVX1 U3375 ( .A(n2734), .Y(n2644) );
  OAI2BB1X1 U3376 ( .A0N(n2734), .A1N(n2660), .B0(n2661), .Y(n2642) );
  XOR3X2 U3377 ( .A(\U3/temp10t[1] ), .B(n2639), .C(\U3/temp12[1] ), .Y(n2655)
         );
  NAND2X1 U3378 ( .A(n2735), .B(n2734), .Y(n2646) );
  XNOR3X2 U3379 ( .A(\U3/temp10t[4] ), .B(\U3/temp10t[3] ), .C(n2636), .Y(
        n2734) );
  XNOR3X2 U3380 ( .A(\U3/temp10t[5] ), .B(n2635), .C(n2634), .Y(n2730) );
  NAND2X1 U3381 ( .A(n2794), .B(n2735), .Y(n2650) );
  XNOR3X2 U3382 ( .A(\U3/temp10t[6] ), .B(\U3/temp10t[5] ), .C(n2633), .Y(
        n2735) );
  OAI21XL U3383 ( .A0(x6[8]), .A1(x1[8]), .B0(n1209), .Y(n1208) );
  NAND2BX1 U3384 ( .AN(\U2/Ytt[10] ), .B(n1254), .Y(\intadd_44/A[7] ) );
  NAND2BX1 U3385 ( .AN(n1302), .B(n2140), .Y(n2449) );
  INVX1 U3386 ( .A(n1316), .Y(n2273) );
  NAND2BX1 U3387 ( .AN(n691), .B(n690), .Y(n2487) );
  OR2X2 U3388 ( .A(n1515), .B(n690), .Y(n2486) );
  XOR3X2 U3389 ( .A(n2694), .B(n2773), .C(n2693), .Y(n2721) );
  XNOR3X2 U3390 ( .A(n2142), .B(n2720), .C(n2213), .Y(n2776) );
  XNOR3X2 U3391 ( .A(n2136), .B(n2813), .C(n2718), .Y(n2291) );
  XNOR3X2 U3392 ( .A(n2144), .B(\U3/temp9t[5] ), .C(n2690), .Y(n2692) );
  XNOR3X2 U3393 ( .A(\U3/temp11[1] ), .B(\U3/temp9t[1] ), .C(n2669), .Y(n2670)
         );
  XNOR3X2 U3394 ( .A(n2144), .B(\U3/temp9t[3] ), .C(n2671), .Y(n2689) );
  XNOR3X2 U3395 ( .A(\U3/temp9t[8] ), .B(n2606), .C(n2681), .Y(n2202) );
  OR2X2 U3396 ( .A(n2555), .B(n749), .Y(n2259) );
  INVX1 U3397 ( .A(n1477), .Y(n2412) );
  AOI22X1 U3398 ( .A0(n1019), .A1(n974), .B0(\U4/U5/temp[11] ), .B1(
        \U4/U5/temp[7] ), .Y(n2267) );
  INVX1 U3399 ( .A(n1483), .Y(n2289) );
  AOI22X1 U3400 ( .A0(n1019), .A1(\U4/U5/temp[5] ), .B0(\U4/U5/temp[11] ), 
        .B1(n1045), .Y(n2185) );
  AOI21X1 U3401 ( .A0(n1352), .A1(n989), .B0(n992), .Y(\U5/Xt[11] ) );
  NAND2X1 U3402 ( .A(n2552), .B(n1877), .Y(n2181) );
  INVX1 U3403 ( .A(n760), .Y(n2594) );
  NAND2X1 U3404 ( .A(n1969), .B(n640), .Y(n2521) );
  NAND2BX1 U3405 ( .AN(n2139), .B(n992), .Y(n2455) );
  INVX1 U3406 ( .A(n1371), .Y(n2249) );
  INVX1 U3407 ( .A(n1374), .Y(n2176) );
  AOI21X1 U3408 ( .A0(n1409), .A1(n977), .B0(n980), .Y(\U4/Yt[11] ) );
  NAND2BX1 U3409 ( .AN(n2138), .B(n980), .Y(n2503) );
  INVX1 U3410 ( .A(n1425), .Y(n2424) );
  INVX1 U3411 ( .A(n1431), .Y(n2361) );
  AOI22X1 U3412 ( .A0(n1020), .A1(\U4/U6/temp[5] ), .B0(\U4/U6/temp[11] ), 
        .B1(n1048), .Y(n2282) );
  NAND2X1 U3413 ( .A(n2543), .B(n1067), .Y(n2351) );
  NAND2X1 U3414 ( .A(n2543), .B(n984), .Y(n2350) );
  NAND2X1 U3415 ( .A(n984), .B(n1067), .Y(n2352) );
  INVX1 U3416 ( .A(n1654), .Y(n2446) );
  INVX1 U3417 ( .A(n1662), .Y(n2317) );
  AOI2BB2X1 U3418 ( .B0(n2561), .B1(n1676), .A0N(n2561), .A1N(n1676), .Y(n1674) );
  XNOR3X2 U3419 ( .A(n2144), .B(\U3/temp9t[9] ), .C(n2679), .Y(n2697) );
  INVX1 U3420 ( .A(n1806), .Y(n2581) );
  XNOR3X2 U3421 ( .A(n2211), .B(n2144), .C(n2683), .Y(n2210) );
  AOI2BB2X1 U3422 ( .B0(n2566), .B1(n1680), .A0N(n2566), .A1N(n1680), .Y(n1678) );
  AOI31X4 U3423 ( .A0(\U4/U5/temp[6] ), .A1(\U4/U5/temp[7] ), .A2(n1493), .B0(
        n1019), .Y(n1463) );
  AOI31X4 U3424 ( .A0(\U4/U6/temp[6] ), .A1(\U4/U6/temp[7] ), .A2(n1441), .B0(
        n1020), .Y(n1411) );
  AOI31X4 U3425 ( .A0(\U5/U5/temp[6] ), .A1(\U5/U5/temp[7] ), .A2(n1384), .B0(
        n1021), .Y(n1354) );
  AOI31X4 U3426 ( .A0(\U5/U6/temp[6] ), .A1(\U5/U6/temp[7] ), .A2(n1332), .B0(
        n1022), .Y(n1302) );
endmodule

